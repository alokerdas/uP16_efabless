magic
tech sky130B
magscale 1 2
timestamp 1659466138
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 404998 700544 405004 700596
rect 405056 700584 405062 700596
rect 413646 700584 413652 700596
rect 405056 700556 413652 700584
rect 405056 700544 405062 700556
rect 413646 700544 413652 700556
rect 413704 700544 413710 700596
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 182818 700516 182824 700528
rect 154172 700488 182824 700516
rect 154172 700476 154178 700488
rect 182818 700476 182824 700488
rect 182876 700476 182882 700528
rect 296070 700476 296076 700528
rect 296128 700516 296134 700528
rect 300118 700516 300124 700528
rect 296128 700488 300124 700516
rect 296128 700476 296134 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 409138 700476 409144 700528
rect 409196 700516 409202 700528
rect 429838 700516 429844 700528
rect 409196 700488 429844 700516
rect 409196 700476 409202 700488
rect 429838 700476 429844 700488
rect 429896 700476 429902 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 178678 700448 178684 700460
rect 137888 700420 178684 700448
rect 137888 700408 137894 700420
rect 178678 700408 178684 700420
rect 178736 700408 178742 700460
rect 188890 700408 188896 700460
rect 188948 700448 188954 700460
rect 202782 700448 202788 700460
rect 188948 700420 202788 700448
rect 188948 700408 188954 700420
rect 202782 700408 202788 700420
rect 202840 700408 202846 700460
rect 293218 700408 293224 700460
rect 293276 700448 293282 700460
rect 332502 700448 332508 700460
rect 293276 700420 332508 700448
rect 293276 700408 293282 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 403618 700408 403624 700460
rect 403676 700448 403682 700460
rect 462314 700448 462320 700460
rect 403676 700420 462320 700448
rect 403676 700408 403682 700420
rect 462314 700408 462320 700420
rect 462372 700408 462378 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 174538 700380 174544 700392
rect 105504 700352 174544 700380
rect 105504 700340 105510 700352
rect 174538 700340 174544 700352
rect 174596 700340 174602 700392
rect 188982 700340 188988 700392
rect 189040 700380 189046 700392
rect 218974 700380 218980 700392
rect 189040 700352 218980 700380
rect 189040 700340 189046 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 291838 700340 291844 700392
rect 291896 700380 291902 700392
rect 348786 700380 348792 700392
rect 291896 700352 348792 700380
rect 291896 700340 291902 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 399478 700340 399484 700392
rect 399536 700380 399542 700392
rect 478506 700380 478512 700392
rect 399536 700352 478512 700380
rect 399536 700340 399542 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 184198 700312 184204 700324
rect 89220 700284 184204 700312
rect 89220 700272 89226 700284
rect 184198 700272 184204 700284
rect 184256 700272 184262 700324
rect 188798 700272 188804 700324
rect 188856 700312 188862 700324
rect 235166 700312 235172 700324
rect 188856 700284 235172 700312
rect 188856 700272 188862 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 283006 700312 283012 700324
rect 267700 700284 283012 700312
rect 267700 700272 267706 700284
rect 283006 700272 283012 700284
rect 283064 700272 283070 700324
rect 295978 700272 295984 700324
rect 296036 700312 296042 700324
rect 364978 700312 364984 700324
rect 296036 700284 364984 700312
rect 296036 700272 296042 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 406378 700272 406384 700324
rect 406436 700312 406442 700324
rect 494790 700312 494796 700324
rect 406436 700284 494796 700312
rect 406436 700272 406442 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 509878 700272 509884 700324
rect 509936 700312 509942 700324
rect 559650 700312 559656 700324
rect 509936 700284 559656 700312
rect 509936 700272 509942 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171778 699700 171784 699712
rect 170364 699672 171784 699700
rect 170364 699660 170370 699672
rect 171778 699660 171784 699672
rect 171836 699660 171842 699712
rect 395338 699660 395344 699712
rect 395396 699700 395402 699712
rect 397454 699700 397460 699712
rect 395396 699672 397460 699700
rect 395396 699660 395402 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 286318 696940 286324 696992
rect 286376 696980 286382 696992
rect 580166 696980 580172 696992
rect 286376 696952 580172 696980
rect 286376 696940 286382 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 508498 670692 508504 670744
rect 508556 670732 508562 670744
rect 580166 670732 580172 670744
rect 508556 670704 580172 670732
rect 508556 670692 508562 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 512638 643084 512644 643136
rect 512696 643124 512702 643136
rect 580166 643124 580172 643136
rect 512696 643096 580172 643124
rect 512696 643084 512702 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 501598 630640 501604 630692
rect 501656 630680 501662 630692
rect 579982 630680 579988 630692
rect 501656 630652 579988 630680
rect 501656 630640 501662 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 504358 616836 504364 616888
rect 504416 616876 504422 616888
rect 580166 616876 580172 616888
rect 504416 616848 580172 616876
rect 504416 616836 504422 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 297358 600108 297364 600160
rect 297416 600148 297422 600160
rect 297910 600148 297916 600160
rect 297416 600120 297916 600148
rect 297416 600108 297422 600120
rect 297910 600108 297916 600120
rect 297968 600108 297974 600160
rect 78122 599972 78128 600024
rect 78180 600012 78186 600024
rect 187234 600012 187240 600024
rect 78180 599984 187240 600012
rect 78180 599972 78186 599984
rect 187234 599972 187240 599984
rect 187292 599972 187298 600024
rect 297928 600012 297956 600108
rect 408126 600012 408132 600024
rect 297928 599984 408132 600012
rect 408126 599972 408132 599984
rect 408184 599972 408190 600024
rect 78030 599904 78036 599956
rect 78088 599944 78094 599956
rect 187142 599944 187148 599956
rect 78088 599916 187148 599944
rect 78088 599904 78094 599916
rect 187142 599904 187148 599916
rect 187200 599904 187206 599956
rect 78582 599836 78588 599888
rect 78640 599876 78646 599888
rect 187326 599876 187332 599888
rect 78640 599848 187332 599876
rect 78640 599836 78646 599848
rect 187326 599836 187332 599848
rect 187384 599836 187390 599888
rect 78214 599768 78220 599820
rect 78272 599808 78278 599820
rect 186866 599808 186872 599820
rect 78272 599780 186872 599808
rect 78272 599768 78278 599780
rect 186866 599768 186872 599780
rect 186924 599768 186930 599820
rect 78490 599700 78496 599752
rect 78548 599740 78554 599752
rect 186958 599740 186964 599752
rect 78548 599712 186964 599740
rect 78548 599700 78554 599712
rect 186958 599700 186964 599712
rect 187016 599700 187022 599752
rect 78398 599632 78404 599684
rect 78456 599672 78462 599684
rect 187050 599672 187056 599684
rect 78456 599644 187056 599672
rect 78456 599632 78462 599644
rect 187050 599632 187056 599644
rect 187108 599632 187114 599684
rect 297450 598884 297456 598936
rect 297508 598924 297514 598936
rect 408218 598924 408224 598936
rect 297508 598896 408224 598924
rect 297508 598884 297514 598896
rect 408218 598884 408224 598896
rect 408276 598884 408282 598936
rect 298002 598816 298008 598868
rect 298060 598856 298066 598868
rect 407942 598856 407948 598868
rect 298060 598828 407948 598856
rect 298060 598816 298066 598828
rect 407942 598816 407948 598828
rect 408000 598816 408006 598868
rect 297542 598748 297548 598800
rect 297600 598788 297606 598800
rect 407574 598788 407580 598800
rect 297600 598760 407580 598788
rect 297600 598748 297606 598760
rect 407574 598748 407580 598760
rect 407632 598748 407638 598800
rect 297266 598544 297272 598596
rect 297324 598584 297330 598596
rect 298002 598584 298008 598596
rect 297324 598556 298008 598584
rect 297324 598544 297330 598556
rect 298002 598544 298008 598556
rect 298060 598544 298066 598596
rect 280982 597320 280988 597372
rect 281040 597360 281046 597372
rect 335354 597360 335360 597372
rect 281040 597332 335360 597360
rect 281040 597320 281046 597332
rect 335354 597320 335360 597332
rect 335412 597320 335418 597372
rect 102870 597252 102876 597304
rect 102928 597292 102934 597304
rect 212350 597292 212356 597304
rect 102928 597264 212356 597292
rect 102928 597252 102934 597264
rect 212350 597252 212356 597264
rect 212408 597252 212414 597304
rect 319990 597252 319996 597304
rect 320048 597292 320054 597304
rect 427814 597292 427820 597304
rect 320048 597264 427820 597292
rect 320048 597252 320054 597264
rect 427814 597252 427820 597264
rect 427872 597252 427878 597304
rect 104802 597184 104808 597236
rect 104860 597224 104866 597236
rect 214834 597224 214840 597236
rect 104860 597196 214840 597224
rect 104860 597184 104866 597196
rect 214834 597184 214840 597196
rect 214892 597184 214898 597236
rect 326154 597184 326160 597236
rect 326212 597224 326218 597236
rect 434714 597224 434720 597236
rect 326212 597196 434720 597224
rect 326212 597184 326218 597196
rect 434714 597184 434720 597196
rect 434772 597184 434778 597236
rect 100662 597116 100668 597168
rect 100720 597156 100726 597168
rect 209958 597156 209964 597168
rect 100720 597128 209964 597156
rect 100720 597116 100726 597128
rect 209958 597116 209964 597128
rect 210016 597156 210022 597168
rect 211062 597156 211068 597168
rect 210016 597128 211068 597156
rect 210016 597116 210022 597128
rect 211062 597116 211068 597128
rect 211120 597116 211126 597168
rect 318702 597116 318708 597168
rect 318760 597156 318766 597168
rect 426434 597156 426440 597168
rect 318760 597128 426440 597156
rect 318760 597116 318766 597128
rect 426434 597116 426440 597128
rect 426492 597116 426498 597168
rect 99282 597048 99288 597100
rect 99340 597088 99346 597100
rect 208946 597088 208952 597100
rect 99340 597060 208952 597088
rect 99340 597048 99346 597060
rect 208946 597048 208952 597060
rect 209004 597048 209010 597100
rect 324406 597048 324412 597100
rect 324464 597088 324470 597100
rect 434714 597088 434720 597100
rect 324464 597060 434720 597088
rect 324464 597048 324470 597060
rect 434714 597048 434720 597060
rect 434772 597048 434778 597100
rect 102042 596980 102048 597032
rect 102100 597020 102106 597032
rect 211154 597020 211160 597032
rect 102100 596992 211160 597020
rect 102100 596980 102106 596992
rect 211154 596980 211160 596992
rect 211212 597020 211218 597032
rect 212442 597020 212448 597032
rect 211212 596992 212448 597020
rect 211212 596980 211218 596992
rect 212442 596980 212448 596992
rect 212500 596980 212506 597032
rect 213822 596980 213828 597032
rect 213880 597020 213886 597032
rect 284570 597020 284576 597032
rect 213880 596992 284576 597020
rect 213880 596980 213886 596992
rect 284570 596980 284576 596992
rect 284628 596980 284634 597032
rect 322934 596980 322940 597032
rect 322992 597020 322998 597032
rect 433334 597020 433340 597032
rect 322992 596992 433340 597020
rect 322992 596980 322998 596992
rect 433334 596980 433340 596992
rect 433392 596980 433398 597032
rect 106182 596912 106188 596964
rect 106240 596952 106246 596964
rect 215754 596952 215760 596964
rect 106240 596924 215760 596952
rect 106240 596912 106246 596924
rect 215754 596912 215760 596924
rect 215812 596952 215818 596964
rect 284386 596952 284392 596964
rect 215812 596924 284392 596952
rect 215812 596912 215818 596924
rect 284386 596912 284392 596924
rect 284444 596912 284450 596964
rect 320910 596912 320916 596964
rect 320968 596952 320974 596964
rect 430574 596952 430580 596964
rect 320968 596924 430580 596952
rect 320968 596912 320974 596924
rect 430574 596912 430580 596924
rect 430632 596912 430638 596964
rect 103422 596844 103428 596896
rect 103480 596884 103486 596896
rect 213822 596884 213828 596896
rect 103480 596856 213828 596884
rect 103480 596844 103486 596856
rect 213822 596844 213828 596856
rect 213880 596844 213886 596896
rect 214834 596844 214840 596896
rect 214892 596884 214898 596896
rect 284478 596884 284484 596896
rect 214892 596856 284484 596884
rect 214892 596844 214898 596856
rect 284478 596844 284484 596856
rect 284536 596844 284542 596896
rect 299290 596844 299296 596896
rect 299348 596884 299354 596896
rect 313274 596884 313280 596896
rect 299348 596856 313280 596884
rect 299348 596844 299354 596856
rect 313274 596844 313280 596856
rect 313332 596844 313338 596896
rect 429194 596884 429200 596896
rect 320560 596856 429200 596884
rect 97902 596776 97908 596828
rect 97960 596816 97966 596828
rect 207842 596816 207848 596828
rect 97960 596788 207848 596816
rect 97960 596776 97966 596788
rect 207842 596776 207848 596788
rect 207900 596776 207906 596828
rect 212442 596776 212448 596828
rect 212500 596816 212506 596828
rect 283190 596816 283196 596828
rect 212500 596788 283196 596816
rect 212500 596776 212506 596788
rect 283190 596776 283196 596788
rect 283248 596776 283254 596828
rect 299198 596776 299204 596828
rect 299256 596816 299262 596828
rect 314654 596816 314660 596828
rect 299256 596788 314660 596816
rect 299256 596776 299262 596788
rect 314654 596776 314660 596788
rect 314712 596776 314718 596828
rect 281074 596708 281080 596760
rect 281132 596748 281138 596760
rect 317690 596748 317696 596760
rect 281132 596720 317696 596748
rect 281132 596708 281138 596720
rect 317690 596708 317696 596720
rect 317748 596748 317754 596760
rect 318702 596748 318708 596760
rect 317748 596720 318708 596748
rect 317748 596708 317754 596720
rect 318702 596708 318708 596720
rect 318760 596708 318766 596760
rect 283098 596640 283104 596692
rect 283156 596680 283162 596692
rect 320082 596680 320088 596692
rect 283156 596652 320088 596680
rect 283156 596640 283162 596652
rect 320082 596640 320088 596652
rect 320140 596680 320146 596692
rect 320560 596680 320588 596856
rect 429194 596844 429200 596856
rect 429252 596844 429258 596896
rect 431954 596816 431960 596828
rect 320140 596652 320588 596680
rect 325666 596788 431960 596816
rect 320140 596640 320146 596652
rect 283190 596572 283196 596624
rect 283248 596612 283254 596624
rect 320910 596612 320916 596624
rect 283248 596584 320916 596612
rect 283248 596572 283254 596584
rect 320910 596572 320916 596584
rect 320968 596572 320974 596624
rect 140682 596504 140688 596556
rect 140740 596544 140746 596556
rect 172146 596544 172152 596556
rect 140740 596516 172152 596544
rect 140740 596504 140746 596516
rect 172146 596504 172152 596516
rect 172204 596504 172210 596556
rect 284294 596504 284300 596556
rect 284352 596544 284358 596556
rect 322198 596544 322204 596556
rect 284352 596516 322204 596544
rect 284352 596504 284358 596516
rect 322198 596504 322204 596516
rect 322256 596544 322262 596556
rect 325666 596544 325694 596788
rect 431954 596776 431960 596788
rect 432012 596776 432018 596828
rect 322256 596516 325694 596544
rect 322256 596504 322262 596516
rect 407942 596504 407948 596556
rect 408000 596544 408006 596556
rect 422570 596544 422576 596556
rect 408000 596516 422576 596544
rect 408000 596504 408006 596516
rect 422570 596504 422576 596516
rect 422628 596504 422634 596556
rect 136542 596436 136548 596488
rect 136600 596476 136606 596488
rect 173342 596476 173348 596488
rect 136600 596448 173348 596476
rect 136600 596436 136606 596448
rect 173342 596436 173348 596448
rect 173400 596436 173406 596488
rect 281534 596436 281540 596488
rect 281592 596476 281598 596488
rect 319990 596476 319996 596488
rect 281592 596448 319996 596476
rect 281592 596436 281598 596448
rect 319990 596436 319996 596448
rect 320048 596436 320054 596488
rect 408126 596436 408132 596488
rect 408184 596476 408190 596488
rect 423674 596476 423680 596488
rect 408184 596448 423680 596476
rect 408184 596436 408190 596448
rect 423674 596436 423680 596448
rect 423732 596436 423738 596488
rect 131022 596368 131028 596420
rect 131080 596408 131086 596420
rect 171870 596408 171876 596420
rect 131080 596380 171876 596408
rect 131080 596368 131086 596380
rect 171870 596368 171876 596380
rect 171928 596368 171934 596420
rect 212350 596368 212356 596420
rect 212408 596408 212414 596420
rect 284294 596408 284300 596420
rect 212408 596380 284300 596408
rect 212408 596368 212414 596380
rect 284294 596368 284300 596380
rect 284352 596368 284358 596420
rect 284570 596368 284576 596420
rect 284628 596408 284634 596420
rect 322934 596408 322940 596420
rect 284628 596380 322940 596408
rect 284628 596368 284634 596380
rect 322934 596368 322940 596380
rect 322992 596368 322998 596420
rect 408218 596368 408224 596420
rect 408276 596408 408282 596420
rect 425054 596408 425060 596420
rect 408276 596380 425060 596408
rect 408276 596368 408282 596380
rect 425054 596368 425060 596380
rect 425112 596368 425118 596420
rect 79778 596300 79784 596352
rect 79836 596340 79842 596352
rect 92474 596340 92480 596352
rect 79836 596312 92480 596340
rect 79836 596300 79842 596312
rect 92474 596300 92480 596312
rect 92532 596300 92538 596352
rect 126882 596300 126888 596352
rect 126940 596340 126946 596352
rect 173250 596340 173256 596352
rect 126940 596312 173256 596340
rect 126940 596300 126946 596312
rect 173250 596300 173256 596312
rect 173308 596300 173314 596352
rect 188614 596300 188620 596352
rect 188672 596340 188678 596352
rect 202874 596340 202880 596352
rect 188672 596312 202880 596340
rect 188672 596300 188678 596312
rect 202874 596300 202880 596312
rect 202932 596300 202938 596352
rect 208946 596300 208952 596352
rect 209004 596340 209010 596352
rect 281534 596340 281540 596352
rect 209004 596312 281540 596340
rect 209004 596300 209010 596312
rect 281534 596300 281540 596312
rect 281592 596300 281598 596352
rect 284478 596300 284484 596352
rect 284536 596340 284542 596352
rect 324406 596340 324412 596352
rect 284536 596312 324412 596340
rect 284536 596300 284542 596312
rect 324406 596300 324412 596312
rect 324464 596300 324470 596352
rect 406470 596300 406476 596352
rect 406528 596340 406534 596352
rect 434714 596340 434720 596352
rect 406528 596312 434720 596340
rect 406528 596300 406534 596312
rect 434714 596300 434720 596312
rect 434772 596300 434778 596352
rect 79962 596232 79968 596284
rect 80020 596272 80026 596284
rect 94038 596272 94044 596284
rect 80020 596244 94044 596272
rect 80020 596232 80026 596244
rect 94038 596232 94044 596244
rect 94096 596232 94102 596284
rect 121362 596232 121368 596284
rect 121420 596272 121426 596284
rect 171962 596272 171968 596284
rect 121420 596244 171968 596272
rect 121420 596232 121426 596244
rect 171962 596232 171968 596244
rect 172020 596232 172026 596284
rect 188706 596232 188712 596284
rect 188764 596272 188770 596284
rect 204346 596272 204352 596284
rect 188764 596244 204352 596272
rect 188764 596232 188770 596244
rect 204346 596232 204352 596244
rect 204404 596232 204410 596284
rect 211062 596232 211068 596284
rect 211120 596272 211126 596284
rect 283098 596272 283104 596284
rect 211120 596244 283104 596272
rect 211120 596232 211126 596244
rect 283098 596232 283104 596244
rect 283156 596232 283162 596284
rect 284386 596232 284392 596284
rect 284444 596272 284450 596284
rect 326154 596272 326160 596284
rect 284444 596244 326160 596272
rect 284444 596232 284450 596244
rect 326154 596232 326160 596244
rect 326212 596232 326218 596284
rect 409414 596232 409420 596284
rect 409472 596272 409478 596284
rect 444374 596272 444380 596284
rect 409472 596244 444380 596272
rect 409472 596232 409478 596244
rect 444374 596232 444380 596244
rect 444432 596232 444438 596284
rect 79870 596164 79876 596216
rect 79928 596204 79934 596216
rect 95234 596204 95240 596216
rect 79928 596176 95240 596204
rect 79928 596164 79934 596176
rect 95234 596164 95240 596176
rect 95292 596164 95298 596216
rect 115842 596164 115848 596216
rect 115900 596204 115906 596216
rect 172054 596204 172060 596216
rect 115900 596176 172060 596204
rect 115900 596164 115906 596176
rect 172054 596164 172060 596176
rect 172112 596164 172118 596216
rect 188522 596164 188528 596216
rect 188580 596204 188586 596216
rect 204254 596204 204260 596216
rect 188580 596176 204260 596204
rect 188580 596164 188586 596176
rect 204254 596164 204260 596176
rect 204312 596164 204318 596216
rect 207842 596164 207848 596216
rect 207900 596204 207906 596216
rect 281074 596204 281080 596216
rect 207900 596176 281080 596204
rect 207900 596164 207906 596176
rect 281074 596164 281080 596176
rect 281132 596164 281138 596216
rect 299382 596164 299388 596216
rect 299440 596204 299446 596216
rect 311894 596204 311900 596216
rect 299440 596176 311900 596204
rect 299440 596164 299446 596176
rect 311894 596164 311900 596176
rect 311952 596164 311958 596216
rect 409230 596164 409236 596216
rect 409288 596204 409294 596216
rect 455414 596204 455420 596216
rect 409288 596176 455420 596204
rect 409288 596164 409294 596176
rect 455414 596164 455420 596176
rect 455472 596164 455478 596216
rect 282178 592628 282184 592680
rect 282236 592668 282242 592680
rect 440234 592668 440240 592680
rect 282236 592640 440240 592668
rect 282236 592628 282242 592640
rect 440234 592628 440240 592640
rect 440292 592628 440298 592680
rect 285030 590656 285036 590708
rect 285088 590696 285094 590708
rect 580166 590696 580172 590708
rect 285088 590668 580172 590696
rect 285088 590656 285094 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 289078 589908 289084 589960
rect 289136 589948 289142 589960
rect 329834 589948 329840 589960
rect 289136 589920 329840 589948
rect 289136 589908 289142 589920
rect 329834 589908 329840 589920
rect 329892 589908 329898 589960
rect 284938 588548 284944 588600
rect 284996 588588 285002 588600
rect 339494 588588 339500 588600
rect 284996 588560 339500 588588
rect 284996 588548 285002 588560
rect 339494 588548 339500 588560
rect 339552 588548 339558 588600
rect 287698 587188 287704 587240
rect 287756 587228 287762 587240
rect 324314 587228 324320 587240
rect 287756 587200 324320 587228
rect 287756 587188 287762 587200
rect 324314 587188 324320 587200
rect 324372 587188 324378 587240
rect 282270 587120 282276 587172
rect 282328 587160 282334 587172
rect 449894 587160 449900 587172
rect 282328 587132 449900 587160
rect 282328 587120 282334 587132
rect 449894 587120 449900 587132
rect 449952 587120 449958 587172
rect 286410 585828 286416 585880
rect 286468 585868 286474 585880
rect 360194 585868 360200 585880
rect 286468 585840 360200 585868
rect 286468 585828 286474 585840
rect 360194 585828 360200 585840
rect 360252 585828 360258 585880
rect 297174 585760 297180 585812
rect 297232 585800 297238 585812
rect 407666 585800 407672 585812
rect 297232 585772 407672 585800
rect 297232 585760 297238 585772
rect 407666 585760 407672 585772
rect 407724 585760 407730 585812
rect 78306 584400 78312 584452
rect 78364 584440 78370 584452
rect 186774 584440 186780 584452
rect 78364 584412 186780 584440
rect 78364 584400 78370 584412
rect 186774 584400 186780 584412
rect 186832 584400 186838 584452
rect 298738 584400 298744 584452
rect 298796 584440 298802 584452
rect 354674 584440 354680 584452
rect 298796 584412 354680 584440
rect 298796 584400 298802 584412
rect 354674 584400 354680 584412
rect 354732 584400 354738 584452
rect 291930 582972 291936 583024
rect 291988 583012 291994 583024
rect 349154 583012 349160 583024
rect 291988 582984 349160 583012
rect 291988 582972 291994 582984
rect 349154 582972 349160 582984
rect 349212 582972 349218 583024
rect 111702 581612 111708 581664
rect 111760 581652 111766 581664
rect 188338 581652 188344 581664
rect 111760 581624 188344 581652
rect 111760 581612 111766 581624
rect 188338 581612 188344 581624
rect 188396 581612 188402 581664
rect 226242 581612 226248 581664
rect 226300 581652 226306 581664
rect 281626 581652 281632 581664
rect 226300 581624 281632 581652
rect 226300 581612 226306 581624
rect 281626 581612 281632 581624
rect 281684 581612 281690 581664
rect 289170 581612 289176 581664
rect 289228 581652 289234 581664
rect 345014 581652 345020 581664
rect 289228 581624 345020 581652
rect 289228 581612 289234 581624
rect 345014 581612 345020 581624
rect 345072 581612 345078 581664
rect 251082 580524 251088 580576
rect 251140 580564 251146 580576
rect 281718 580564 281724 580576
rect 251140 580536 281724 580564
rect 251140 580524 251146 580536
rect 281718 580524 281724 580536
rect 281776 580524 281782 580576
rect 245562 580456 245568 580508
rect 245620 580496 245626 580508
rect 281810 580496 281816 580508
rect 245620 580468 281816 580496
rect 245620 580456 245626 580468
rect 281810 580456 281816 580468
rect 281868 580456 281874 580508
rect 241422 580388 241428 580440
rect 241480 580428 241486 580440
rect 282086 580428 282092 580440
rect 241480 580400 282092 580428
rect 241480 580388 241486 580400
rect 282086 580388 282092 580400
rect 282144 580388 282150 580440
rect 189994 580320 190000 580372
rect 190052 580360 190058 580372
rect 215294 580360 215300 580372
rect 190052 580332 215300 580360
rect 190052 580320 190058 580332
rect 215294 580320 215300 580332
rect 215352 580320 215358 580372
rect 235902 580320 235908 580372
rect 235960 580360 235966 580372
rect 281902 580360 281908 580372
rect 235960 580332 281908 580360
rect 235960 580320 235966 580332
rect 281902 580320 281908 580332
rect 281960 580320 281966 580372
rect 189902 580252 189908 580304
rect 189960 580292 189966 580304
rect 219434 580292 219440 580304
rect 189960 580264 219440 580292
rect 189960 580252 189966 580264
rect 219434 580252 219440 580264
rect 219492 580252 219498 580304
rect 231762 580252 231768 580304
rect 231820 580292 231826 580304
rect 281994 580292 282000 580304
rect 231820 580264 282000 580292
rect 231820 580252 231826 580264
rect 281994 580252 282000 580264
rect 282052 580252 282058 580304
rect 282362 580252 282368 580304
rect 282420 580292 282426 580304
rect 459554 580292 459560 580304
rect 282420 580264 459560 580292
rect 282420 580252 282426 580264
rect 459554 580252 459560 580264
rect 459612 580252 459618 580304
rect 516778 576852 516784 576904
rect 516836 576892 516842 576904
rect 580166 576892 580172 576904
rect 516836 576864 580172 576892
rect 516836 576852 516842 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3326 565836 3332 565888
rect 3384 565876 3390 565888
rect 32398 565876 32404 565888
rect 3384 565848 32404 565876
rect 3384 565836 3390 565848
rect 32398 565836 32404 565848
rect 32456 565836 32462 565888
rect 507118 563048 507124 563100
rect 507176 563088 507182 563100
rect 580166 563088 580172 563100
rect 507176 563060 580172 563088
rect 507176 563048 507182 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3142 553392 3148 553444
rect 3200 553432 3206 553444
rect 22738 553432 22744 553444
rect 3200 553404 22744 553432
rect 3200 553392 3206 553404
rect 22738 553392 22744 553404
rect 22796 553392 22802 553444
rect 511258 536800 511264 536852
rect 511316 536840 511322 536852
rect 579890 536840 579896 536852
rect 511316 536812 579896 536840
rect 511316 536800 511322 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 14458 527184 14464 527196
rect 3384 527156 14464 527184
rect 3384 527144 3390 527156
rect 14458 527144 14464 527156
rect 14516 527144 14522 527196
rect 293862 526736 293868 526788
rect 293920 526776 293926 526788
rect 297266 526776 297272 526788
rect 293920 526748 297272 526776
rect 293920 526736 293926 526748
rect 297266 526736 297272 526748
rect 297324 526776 297330 526788
rect 298002 526776 298008 526788
rect 297324 526748 298008 526776
rect 297324 526736 297330 526748
rect 298002 526736 298008 526748
rect 298060 526736 298066 526788
rect 187326 525784 187332 525836
rect 187384 525824 187390 525836
rect 187694 525824 187700 525836
rect 187384 525796 187700 525824
rect 187384 525784 187390 525796
rect 187694 525784 187700 525796
rect 187752 525784 187758 525836
rect 514018 524424 514024 524476
rect 514076 524464 514082 524476
rect 580166 524464 580172 524476
rect 514076 524436 580172 524464
rect 514076 524424 514082 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 502978 510620 502984 510672
rect 503036 510660 503042 510672
rect 580166 510660 580172 510672
rect 503036 510632 580172 510660
rect 503036 510620 503042 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 10318 501004 10324 501016
rect 3292 500976 10324 501004
rect 3292 500964 3298 500976
rect 10318 500964 10324 500976
rect 10376 500964 10382 501016
rect 287790 498788 287796 498840
rect 287848 498828 287854 498840
rect 296990 498828 296996 498840
rect 287848 498800 296996 498828
rect 287848 498788 287854 498800
rect 296990 498788 296996 498800
rect 297048 498828 297054 498840
rect 297818 498828 297824 498840
rect 297048 498800 297824 498828
rect 297048 498788 297054 498800
rect 297818 498788 297824 498800
rect 297876 498788 297882 498840
rect 187050 493348 187056 493400
rect 187108 493348 187114 493400
rect 187068 493320 187096 493348
rect 187068 493292 187188 493320
rect 186682 493212 186688 493264
rect 186740 493252 186746 493264
rect 187050 493252 187056 493264
rect 186740 493224 187056 493252
rect 186740 493212 186746 493224
rect 187050 493212 187056 493224
rect 187108 493212 187114 493264
rect 186866 493076 186872 493128
rect 186924 493116 186930 493128
rect 187160 493116 187188 493292
rect 186924 493088 187188 493116
rect 186924 493076 186930 493088
rect 78490 489812 78496 489864
rect 78548 489852 78554 489864
rect 187694 489852 187700 489864
rect 78548 489824 187700 489852
rect 78548 489812 78554 489824
rect 187694 489812 187700 489824
rect 187752 489812 187758 489864
rect 297450 489812 297456 489864
rect 297508 489852 297514 489864
rect 297726 489852 297732 489864
rect 297508 489824 297732 489852
rect 297508 489812 297514 489824
rect 297726 489812 297732 489824
rect 297784 489852 297790 489864
rect 407666 489852 407672 489864
rect 297784 489824 407672 489852
rect 297784 489812 297790 489824
rect 407666 489812 407672 489824
rect 407724 489812 407730 489864
rect 77662 489744 77668 489796
rect 77720 489784 77726 489796
rect 187234 489784 187240 489796
rect 77720 489756 187240 489784
rect 77720 489744 77726 489756
rect 187234 489744 187240 489756
rect 187292 489744 187298 489796
rect 78398 489676 78404 489728
rect 78456 489716 78462 489728
rect 187050 489716 187056 489728
rect 78456 489688 187056 489716
rect 78456 489676 78462 489688
rect 187050 489676 187056 489688
rect 187108 489676 187114 489728
rect 78306 489608 78312 489660
rect 78364 489648 78370 489660
rect 187326 489648 187332 489660
rect 78364 489620 187332 489648
rect 78364 489608 78370 489620
rect 187326 489608 187332 489620
rect 187384 489608 187390 489660
rect 78122 489540 78128 489592
rect 78180 489580 78186 489592
rect 186958 489580 186964 489592
rect 78180 489552 186964 489580
rect 78180 489540 78186 489552
rect 186958 489540 186964 489552
rect 187016 489540 187022 489592
rect 77754 489472 77760 489524
rect 77812 489512 77818 489524
rect 186774 489512 186780 489524
rect 77812 489484 186780 489512
rect 77812 489472 77818 489484
rect 186774 489472 186780 489484
rect 186832 489472 186838 489524
rect 78030 489404 78036 489456
rect 78088 489444 78094 489456
rect 186866 489444 186872 489456
rect 78088 489416 186872 489444
rect 78088 489404 78094 489416
rect 186866 489404 186872 489416
rect 186924 489404 186930 489456
rect 78582 489336 78588 489388
rect 78640 489376 78646 489388
rect 187142 489376 187148 489388
rect 78640 489348 187148 489376
rect 78640 489336 78646 489348
rect 187142 489336 187148 489348
rect 187200 489336 187206 489388
rect 173342 489200 173348 489252
rect 173400 489240 173406 489252
rect 253658 489240 253664 489252
rect 173400 489212 253664 489240
rect 173400 489200 173406 489212
rect 253658 489200 253664 489212
rect 253716 489200 253722 489252
rect 218054 489132 218060 489184
rect 218112 489172 218118 489184
rect 404998 489172 405004 489184
rect 218112 489144 405004 489172
rect 218112 489132 218118 489144
rect 404998 489132 405004 489144
rect 405056 489132 405062 489184
rect 186866 488724 186872 488776
rect 186924 488764 186930 488776
rect 187602 488764 187608 488776
rect 186924 488736 187608 488764
rect 186924 488724 186930 488736
rect 187602 488724 187608 488736
rect 187660 488724 187666 488776
rect 187234 488656 187240 488708
rect 187292 488696 187298 488708
rect 187510 488696 187516 488708
rect 187292 488668 187516 488696
rect 187292 488656 187298 488668
rect 187510 488656 187516 488668
rect 187568 488656 187574 488708
rect 187050 488588 187056 488640
rect 187108 488628 187114 488640
rect 187418 488628 187424 488640
rect 187108 488600 187424 488628
rect 187108 488588 187114 488600
rect 187418 488588 187424 488600
rect 187476 488588 187482 488640
rect 186774 488520 186780 488572
rect 186832 488560 186838 488572
rect 187234 488560 187240 488572
rect 186832 488532 187240 488560
rect 186832 488520 186838 488532
rect 187234 488520 187240 488532
rect 187292 488520 187298 488572
rect 79778 488452 79784 488504
rect 79836 488492 79842 488504
rect 92934 488492 92940 488504
rect 79836 488464 92940 488492
rect 79836 488452 79842 488464
rect 92934 488452 92940 488464
rect 92992 488492 92998 488504
rect 188614 488492 188620 488504
rect 92992 488464 188620 488492
rect 92992 488452 92998 488464
rect 188614 488452 188620 488464
rect 188672 488452 188678 488504
rect 297082 488452 297088 488504
rect 297140 488492 297146 488504
rect 297542 488492 297548 488504
rect 297140 488464 297548 488492
rect 297140 488452 297146 488464
rect 297542 488452 297548 488464
rect 297600 488452 297606 488504
rect 297726 488452 297732 488504
rect 297784 488492 297790 488504
rect 298002 488492 298008 488504
rect 297784 488464 298008 488492
rect 297784 488452 297790 488464
rect 298002 488452 298008 488464
rect 298060 488452 298066 488504
rect 408218 488452 408224 488504
rect 408276 488492 408282 488504
rect 425054 488492 425060 488504
rect 408276 488464 425060 488492
rect 408276 488452 408282 488464
rect 425054 488452 425060 488464
rect 425112 488452 425118 488504
rect 79962 488384 79968 488436
rect 80020 488424 80026 488436
rect 94222 488424 94228 488436
rect 80020 488396 94228 488424
rect 80020 488384 80026 488396
rect 94222 488384 94228 488396
rect 94280 488424 94286 488436
rect 188522 488424 188528 488436
rect 94280 488396 188528 488424
rect 94280 488384 94286 488396
rect 188522 488384 188528 488396
rect 188580 488424 188586 488436
rect 204714 488424 204720 488436
rect 188580 488396 204720 488424
rect 188580 488384 188586 488396
rect 204714 488384 204720 488396
rect 204772 488384 204778 488436
rect 292022 488384 292028 488436
rect 292080 488424 292086 488436
rect 297634 488424 297640 488436
rect 292080 488396 297640 488424
rect 292080 488384 292086 488396
rect 297634 488384 297640 488396
rect 297692 488424 297698 488436
rect 407850 488424 407856 488436
rect 297692 488396 407856 488424
rect 297692 488384 297698 488396
rect 407850 488384 407856 488396
rect 407908 488384 407914 488436
rect 408126 488384 408132 488436
rect 408184 488424 408190 488436
rect 423674 488424 423680 488436
rect 408184 488396 423680 488424
rect 408184 488384 408190 488396
rect 423674 488384 423680 488396
rect 423732 488384 423738 488436
rect 79870 488316 79876 488368
rect 79928 488356 79934 488368
rect 95326 488356 95332 488368
rect 79928 488328 95332 488356
rect 79928 488316 79934 488328
rect 95326 488316 95332 488328
rect 95384 488356 95390 488368
rect 95384 488328 180794 488356
rect 95384 488316 95390 488328
rect 180766 488152 180794 488328
rect 298002 488316 298008 488368
rect 298060 488356 298066 488368
rect 407758 488356 407764 488368
rect 298060 488328 407764 488356
rect 298060 488316 298066 488328
rect 407758 488316 407764 488328
rect 407816 488316 407822 488368
rect 407942 488316 407948 488368
rect 408000 488356 408006 488368
rect 422570 488356 422576 488368
rect 408000 488328 422576 488356
rect 408000 488316 408006 488328
rect 422570 488316 422576 488328
rect 422628 488316 422634 488368
rect 298094 488248 298100 488300
rect 298152 488288 298158 488300
rect 299290 488288 299296 488300
rect 298152 488260 299296 488288
rect 298152 488248 298158 488260
rect 299290 488248 299296 488260
rect 299348 488288 299354 488300
rect 314286 488288 314292 488300
rect 299348 488260 314292 488288
rect 299348 488248 299354 488260
rect 314286 488248 314292 488260
rect 314344 488288 314350 488300
rect 408126 488288 408132 488300
rect 314344 488260 408132 488288
rect 314344 488248 314350 488260
rect 408126 488248 408132 488260
rect 408184 488248 408190 488300
rect 188614 488180 188620 488232
rect 188672 488220 188678 488232
rect 202874 488220 202880 488232
rect 188672 488192 202880 488220
rect 188672 488180 188678 488192
rect 202874 488180 202880 488192
rect 202932 488180 202938 488232
rect 299198 488220 299204 488232
rect 292546 488192 299204 488220
rect 188706 488152 188712 488164
rect 180766 488124 188712 488152
rect 188706 488112 188712 488124
rect 188764 488152 188770 488164
rect 204898 488152 204904 488164
rect 188764 488124 204904 488152
rect 188764 488112 188770 488124
rect 204898 488112 204904 488124
rect 204956 488112 204962 488164
rect 188798 488044 188804 488096
rect 188856 488084 188862 488096
rect 220078 488084 220084 488096
rect 188856 488056 220084 488084
rect 188856 488044 188862 488056
rect 220078 488044 220084 488056
rect 220136 488044 220142 488096
rect 105722 487976 105728 488028
rect 105780 488016 105786 488028
rect 215754 488016 215760 488028
rect 105780 487988 215760 488016
rect 105780 487976 105786 487988
rect 215754 487976 215760 487988
rect 215812 487976 215818 488028
rect 230566 487976 230572 488028
rect 230624 488016 230630 488028
rect 287790 488016 287796 488028
rect 230624 487988 287796 488016
rect 230624 487976 230630 487988
rect 287790 487976 287796 487988
rect 287848 487976 287854 488028
rect 104802 487908 104808 487960
rect 104860 487948 104866 487960
rect 214834 487948 214840 487960
rect 104860 487920 214840 487948
rect 104860 487908 104866 487920
rect 214834 487908 214840 487920
rect 214892 487908 214898 487960
rect 219802 487908 219808 487960
rect 219860 487948 219866 487960
rect 283006 487948 283012 487960
rect 219860 487920 283012 487948
rect 219860 487908 219866 487920
rect 283006 487908 283012 487920
rect 283064 487908 283070 487960
rect 103422 487840 103428 487892
rect 103480 487880 103486 487892
rect 213730 487880 213736 487892
rect 103480 487852 213736 487880
rect 103480 487840 103486 487852
rect 213730 487840 213736 487852
rect 213788 487840 213794 487892
rect 232590 487840 232596 487892
rect 232648 487880 232654 487892
rect 292546 487880 292574 488192
rect 299198 488180 299204 488192
rect 299256 488220 299262 488232
rect 315390 488220 315396 488232
rect 299256 488192 315396 488220
rect 299256 488180 299262 488192
rect 315390 488180 315396 488192
rect 315448 488220 315454 488232
rect 408218 488220 408224 488232
rect 315448 488192 408224 488220
rect 315448 488180 315454 488192
rect 408218 488180 408224 488192
rect 408276 488180 408282 488232
rect 297542 488112 297548 488164
rect 297600 488152 297606 488164
rect 408310 488152 408316 488164
rect 297600 488124 408316 488152
rect 297600 488112 297606 488124
rect 408310 488112 408316 488124
rect 408368 488112 408374 488164
rect 232648 487852 292574 487880
rect 232648 487840 232654 487852
rect 101122 487772 101128 487824
rect 101180 487812 101186 487824
rect 211154 487812 211160 487824
rect 101180 487784 211160 487812
rect 101180 487772 101186 487784
rect 211154 487772 211160 487784
rect 211212 487812 211218 487824
rect 212442 487812 212448 487824
rect 211212 487784 212448 487812
rect 211212 487772 211218 487784
rect 212442 487772 212448 487784
rect 212500 487772 212506 487824
rect 232498 487772 232504 487824
rect 232556 487812 232562 487824
rect 298094 487812 298100 487824
rect 232556 487784 298100 487812
rect 232556 487772 232562 487784
rect 298094 487772 298100 487784
rect 298152 487772 298158 487824
rect 312538 487772 312544 487824
rect 312596 487812 312602 487824
rect 312998 487812 313004 487824
rect 312596 487784 313004 487812
rect 312596 487772 312602 487784
rect 312998 487772 313004 487784
rect 313056 487812 313062 487824
rect 407942 487812 407948 487824
rect 313056 487784 407948 487812
rect 313056 487772 313062 487784
rect 407942 487772 407948 487784
rect 408000 487772 408006 487824
rect 326614 487636 326620 487688
rect 326672 487676 326678 487688
rect 434714 487676 434720 487688
rect 326672 487648 434720 487676
rect 326672 487636 326678 487648
rect 434714 487636 434720 487648
rect 434772 487636 434778 487688
rect 319438 487568 319444 487620
rect 319496 487608 319502 487620
rect 427814 487608 427820 487620
rect 319496 487580 427820 487608
rect 319496 487568 319502 487580
rect 427814 487568 427820 487580
rect 427872 487568 427878 487620
rect 318058 487500 318064 487552
rect 318116 487540 318122 487552
rect 426434 487540 426440 487552
rect 318116 487512 426440 487540
rect 318116 487500 318122 487512
rect 426434 487500 426440 487512
rect 426492 487500 426498 487552
rect 97810 487432 97816 487484
rect 97868 487472 97874 487484
rect 207658 487472 207664 487484
rect 97868 487444 207664 487472
rect 97868 487432 97874 487444
rect 207658 487432 207664 487444
rect 207716 487432 207722 487484
rect 214834 487432 214840 487484
rect 214892 487472 214898 487484
rect 228358 487472 228364 487484
rect 214892 487444 228364 487472
rect 214892 487432 214898 487444
rect 228358 487432 228364 487444
rect 228416 487432 228422 487484
rect 319990 487432 319996 487484
rect 320048 487472 320054 487484
rect 429194 487472 429200 487484
rect 320048 487444 429200 487472
rect 320048 487432 320054 487444
rect 429194 487432 429200 487444
rect 429252 487432 429258 487484
rect 102410 487364 102416 487416
rect 102468 487404 102474 487416
rect 212350 487404 212356 487416
rect 102468 487376 212356 487404
rect 102468 487364 102474 487376
rect 212350 487364 212356 487376
rect 212408 487364 212414 487416
rect 212442 487364 212448 487416
rect 212500 487404 212506 487416
rect 226978 487404 226984 487416
rect 212500 487376 226984 487404
rect 212500 487364 212506 487376
rect 226978 487364 226984 487376
rect 227036 487364 227042 487416
rect 322934 487364 322940 487416
rect 322992 487404 322998 487416
rect 433334 487404 433340 487416
rect 322992 487376 433340 487404
rect 322992 487364 322998 487376
rect 433334 487364 433340 487376
rect 433392 487364 433398 487416
rect 98914 487296 98920 487348
rect 98972 487336 98978 487348
rect 208854 487336 208860 487348
rect 98972 487308 208860 487336
rect 98972 487296 98978 487308
rect 208854 487296 208860 487308
rect 208912 487296 208918 487348
rect 213730 487296 213736 487348
rect 213788 487336 213794 487348
rect 229738 487336 229744 487348
rect 213788 487308 229744 487336
rect 213788 487296 213794 487308
rect 229738 487296 229744 487308
rect 229796 487296 229802 487348
rect 324406 487296 324412 487348
rect 324464 487336 324470 487348
rect 434714 487336 434720 487348
rect 324464 487308 434720 487336
rect 324464 487296 324470 487308
rect 434714 487296 434720 487308
rect 434772 487296 434778 487348
rect 204714 487228 204720 487280
rect 204772 487268 204778 487280
rect 222838 487268 222844 487280
rect 204772 487240 222844 487268
rect 204772 487228 204778 487240
rect 222838 487228 222844 487240
rect 222896 487228 222902 487280
rect 322198 487228 322204 487280
rect 322256 487268 322262 487280
rect 432138 487268 432144 487280
rect 322256 487240 432144 487268
rect 322256 487228 322262 487240
rect 432138 487228 432144 487240
rect 432196 487228 432202 487280
rect 100018 487160 100024 487212
rect 100076 487200 100082 487212
rect 210418 487200 210424 487212
rect 100076 487172 210424 487200
rect 100076 487160 100082 487172
rect 210418 487160 210424 487172
rect 210476 487160 210482 487212
rect 215754 487160 215760 487212
rect 215812 487200 215818 487212
rect 244274 487200 244280 487212
rect 215812 487172 244280 487200
rect 215812 487160 215818 487172
rect 244274 487160 244280 487172
rect 244332 487160 244338 487212
rect 320818 487160 320824 487212
rect 320876 487200 320882 487212
rect 430574 487200 430580 487212
rect 320876 487172 430580 487200
rect 320876 487160 320882 487172
rect 430574 487160 430580 487172
rect 430632 487160 430638 487212
rect 436738 487160 436744 487212
rect 436796 487200 436802 487212
rect 465074 487200 465080 487212
rect 436796 487172 465080 487200
rect 436796 487160 436802 487172
rect 465074 487160 465080 487172
rect 465132 487160 465138 487212
rect 299382 487092 299388 487144
rect 299440 487132 299446 487144
rect 311894 487132 311900 487144
rect 299440 487104 311900 487132
rect 299440 487092 299446 487104
rect 311894 487092 311900 487104
rect 311952 487132 311958 487144
rect 312538 487132 312544 487144
rect 311952 487104 312544 487132
rect 311952 487092 311958 487104
rect 312538 487092 312544 487104
rect 312596 487092 312602 487144
rect 246482 486616 246488 486668
rect 246540 486656 246546 486668
rect 249794 486656 249800 486668
rect 246540 486628 249800 486656
rect 246540 486616 246546 486628
rect 249794 486616 249800 486628
rect 249852 486616 249858 486668
rect 208854 486548 208860 486600
rect 208912 486588 208918 486600
rect 238018 486588 238024 486600
rect 208912 486560 238024 486588
rect 208912 486548 208918 486560
rect 238018 486548 238024 486560
rect 238076 486548 238082 486600
rect 244918 486548 244924 486600
rect 244976 486588 244982 486600
rect 324406 486588 324412 486600
rect 244976 486560 324412 486588
rect 244976 486548 244982 486560
rect 324406 486548 324412 486560
rect 324464 486548 324470 486600
rect 187694 486480 187700 486532
rect 187752 486520 187758 486532
rect 235258 486520 235264 486532
rect 187752 486492 235264 486520
rect 187752 486480 187758 486492
rect 235258 486480 235264 486492
rect 235316 486480 235322 486532
rect 248414 486480 248420 486532
rect 248472 486520 248478 486532
rect 409414 486520 409420 486532
rect 248472 486492 409420 486520
rect 248472 486480 248478 486492
rect 409414 486480 409420 486492
rect 409472 486480 409478 486532
rect 216766 486412 216772 486464
rect 216824 486452 216830 486464
rect 542354 486452 542360 486464
rect 216824 486424 542360 486452
rect 216824 486412 216830 486424
rect 542354 486412 542360 486424
rect 542412 486412 542418 486464
rect 243814 485800 243820 485852
rect 243872 485840 243878 485852
rect 244642 485840 244648 485852
rect 243872 485812 244648 485840
rect 243872 485800 243878 485812
rect 244642 485800 244648 485812
rect 244700 485800 244706 485852
rect 239398 485188 239404 485240
rect 239456 485228 239462 485240
rect 319990 485228 319996 485240
rect 239456 485200 319996 485228
rect 239456 485188 239462 485200
rect 319990 485188 319996 485200
rect 320048 485188 320054 485240
rect 172146 485120 172152 485172
rect 172204 485160 172210 485172
rect 254946 485160 254952 485172
rect 172204 485132 254952 485160
rect 172204 485120 172210 485132
rect 254946 485120 254952 485132
rect 255004 485120 255010 485172
rect 253934 485052 253940 485104
rect 253992 485092 253998 485104
rect 409322 485092 409328 485104
rect 253992 485064 409328 485092
rect 253992 485052 253998 485064
rect 409322 485052 409328 485064
rect 409380 485052 409386 485104
rect 221458 484372 221464 484424
rect 221516 484412 221522 484424
rect 580166 484412 580172 484424
rect 221516 484384 580172 484412
rect 221516 484372 221522 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 244274 484304 244280 484356
rect 244332 484344 244338 484356
rect 326614 484344 326620 484356
rect 244332 484316 326620 484344
rect 244332 484304 244338 484316
rect 326614 484304 326620 484316
rect 326672 484304 326678 484356
rect 212350 483692 212356 483744
rect 212408 483732 212414 483744
rect 242158 483732 242164 483744
rect 212408 483704 242164 483732
rect 212408 483692 212414 483704
rect 242158 483692 242164 483704
rect 242216 483692 242222 483744
rect 251174 483692 251180 483744
rect 251232 483732 251238 483744
rect 409230 483732 409236 483744
rect 251232 483704 409236 483732
rect 251232 483692 251238 483704
rect 409230 483692 409236 483704
rect 409288 483692 409294 483744
rect 216950 483624 216956 483676
rect 217008 483664 217014 483676
rect 580258 483664 580264 483676
rect 217008 483636 580264 483664
rect 217008 483624 217014 483636
rect 580258 483624 580264 483636
rect 580316 483624 580322 483676
rect 105814 482332 105820 482384
rect 105872 482372 105878 482384
rect 234614 482372 234620 482384
rect 105872 482344 234620 482372
rect 105872 482332 105878 482344
rect 234614 482332 234620 482344
rect 234672 482332 234678 482384
rect 236086 482332 236092 482384
rect 236144 482372 236150 482384
rect 434714 482372 434720 482384
rect 236144 482344 434720 482372
rect 236144 482332 236150 482344
rect 434714 482332 434720 482344
rect 434772 482332 434778 482384
rect 216674 482264 216680 482316
rect 216732 482304 216738 482316
rect 501598 482304 501604 482316
rect 216732 482276 501604 482304
rect 216732 482264 216738 482276
rect 501598 482264 501604 482276
rect 501656 482264 501662 482316
rect 173250 481108 173256 481160
rect 173308 481148 173314 481160
rect 250806 481148 250812 481160
rect 173308 481120 250812 481148
rect 173308 481108 173314 481120
rect 250806 481108 250812 481120
rect 250864 481108 250870 481160
rect 243538 481040 243544 481092
rect 243596 481080 243602 481092
rect 322934 481080 322940 481092
rect 243596 481052 322940 481080
rect 243596 481040 243602 481052
rect 322934 481040 322940 481052
rect 322992 481040 322998 481092
rect 247862 480972 247868 481024
rect 247920 481012 247926 481024
rect 360194 481012 360200 481024
rect 247920 480984 360200 481012
rect 247920 480972 247926 480984
rect 360194 480972 360200 480984
rect 360252 480972 360258 481024
rect 215294 480904 215300 480956
rect 215352 480944 215358 480956
rect 516778 480944 516784 480956
rect 215352 480916 516784 480944
rect 215352 480904 215358 480916
rect 516778 480904 516784 480916
rect 516836 480904 516842 480956
rect 126882 479680 126888 479732
rect 126940 479720 126946 479732
rect 240870 479720 240876 479732
rect 126940 479692 240876 479720
rect 126940 479680 126946 479692
rect 240870 479680 240876 479692
rect 240928 479680 240934 479732
rect 238846 479612 238852 479664
rect 238904 479652 238910 479664
rect 339494 479652 339500 479664
rect 238904 479624 339500 479652
rect 238904 479612 238910 479624
rect 339494 479612 339500 479624
rect 339552 479612 339558 479664
rect 240778 479544 240784 479596
rect 240836 479584 240842 479596
rect 320818 479584 320824 479596
rect 240836 479556 320824 479584
rect 240836 479544 240842 479556
rect 320818 479544 320824 479556
rect 320876 479544 320882 479596
rect 215478 479476 215484 479528
rect 215536 479516 215542 479528
rect 514018 479516 514024 479528
rect 215536 479488 514024 479516
rect 215536 479476 215542 479488
rect 514018 479476 514024 479488
rect 514076 479476 514082 479528
rect 241422 478932 241428 478984
rect 241480 478972 241486 478984
rect 242250 478972 242256 478984
rect 241480 478944 242256 478972
rect 241480 478932 241486 478944
rect 242250 478932 242256 478944
rect 242308 478932 242314 478984
rect 172054 478252 172060 478304
rect 172112 478292 172118 478304
rect 248506 478292 248512 478304
rect 172112 478264 248512 478292
rect 172112 478252 172118 478264
rect 248506 478252 248512 478264
rect 248564 478252 248570 478304
rect 246574 478184 246580 478236
rect 246632 478224 246638 478236
rect 354674 478224 354680 478236
rect 246632 478196 354680 478224
rect 246632 478184 246638 478196
rect 354674 478184 354680 478196
rect 354732 478184 354738 478236
rect 218238 478116 218244 478168
rect 218296 478156 218302 478168
rect 395338 478156 395344 478168
rect 218296 478128 395344 478156
rect 218296 478116 218302 478128
rect 395338 478116 395344 478128
rect 395396 478116 395402 478168
rect 235258 477436 235264 477488
rect 235316 477476 235322 477488
rect 293310 477476 293316 477488
rect 235316 477448 293316 477476
rect 235316 477436 235322 477448
rect 293310 477436 293316 477448
rect 293368 477436 293374 477488
rect 218146 476824 218152 476876
rect 218204 476864 218210 476876
rect 403618 476864 403624 476876
rect 218204 476836 403624 476864
rect 218204 476824 218210 476836
rect 403618 476824 403624 476836
rect 403676 476824 403682 476876
rect 220722 476756 220728 476808
rect 220780 476796 220786 476808
rect 229830 476796 229836 476808
rect 220780 476768 229836 476796
rect 220780 476756 220786 476768
rect 229830 476756 229836 476768
rect 229888 476756 229894 476808
rect 243630 476756 243636 476808
rect 243688 476796 243694 476808
rect 459554 476796 459560 476808
rect 243688 476768 459560 476796
rect 243688 476756 243694 476768
rect 459554 476756 459560 476768
rect 459612 476756 459618 476808
rect 234798 476076 234804 476128
rect 234856 476116 234862 476128
rect 235258 476116 235264 476128
rect 234856 476088 235264 476116
rect 234856 476076 234862 476088
rect 235258 476076 235264 476088
rect 235316 476076 235322 476128
rect 236546 475464 236552 475516
rect 236604 475504 236610 475516
rect 318058 475504 318064 475516
rect 236604 475476 318064 475504
rect 236604 475464 236610 475476
rect 318058 475464 318064 475476
rect 318116 475464 318122 475516
rect 77938 475396 77944 475448
rect 77996 475436 78002 475448
rect 229922 475436 229928 475448
rect 77996 475408 229928 475436
rect 77996 475396 78002 475408
rect 229922 475396 229928 475408
rect 229980 475396 229986 475448
rect 236270 475396 236276 475448
rect 236328 475436 236334 475448
rect 329834 475436 329840 475448
rect 236328 475408 329840 475436
rect 236328 475396 236334 475408
rect 329834 475396 329840 475408
rect 329892 475396 329898 475448
rect 217134 475328 217140 475380
rect 217192 475368 217198 475380
rect 527174 475368 527180 475380
rect 217192 475340 527180 475368
rect 217192 475328 217198 475340
rect 527174 475328 527180 475340
rect 527232 475328 527238 475380
rect 3234 474716 3240 474768
rect 3292 474756 3298 474768
rect 40678 474756 40684 474768
rect 3292 474728 40684 474756
rect 3292 474716 3298 474728
rect 40678 474716 40684 474728
rect 40736 474716 40742 474768
rect 241606 474648 241612 474700
rect 241664 474688 241670 474700
rect 242158 474688 242164 474700
rect 241664 474660 242164 474688
rect 241664 474648 241670 474660
rect 242158 474648 242164 474660
rect 242216 474688 242222 474700
rect 322198 474688 322204 474700
rect 242216 474660 322204 474688
rect 242216 474648 242222 474660
rect 322198 474648 322204 474660
rect 322256 474648 322262 474700
rect 173158 474104 173164 474156
rect 173216 474144 173222 474156
rect 245654 474144 245660 474156
rect 173216 474116 245660 474144
rect 173216 474104 173222 474116
rect 245654 474104 245660 474116
rect 245712 474104 245718 474156
rect 237742 474036 237748 474088
rect 237800 474076 237806 474088
rect 335354 474076 335360 474088
rect 237800 474048 335360 474076
rect 237800 474036 237806 474048
rect 335354 474036 335360 474048
rect 335412 474036 335418 474088
rect 215662 473968 215668 474020
rect 215720 474008 215726 474020
rect 512638 474008 512644 474020
rect 215720 473980 512644 474008
rect 215720 473968 215726 473980
rect 512638 473968 512644 473980
rect 512696 473968 512702 474020
rect 237558 473288 237564 473340
rect 237616 473328 237622 473340
rect 238018 473328 238024 473340
rect 237616 473300 238024 473328
rect 237616 473288 237622 473300
rect 238018 473288 238024 473300
rect 238076 473328 238082 473340
rect 319438 473328 319444 473340
rect 238076 473300 319444 473328
rect 238076 473288 238082 473300
rect 319438 473288 319444 473300
rect 319496 473288 319502 473340
rect 235902 473016 235908 473068
rect 235960 473056 235966 473068
rect 240962 473056 240968 473068
rect 235960 473028 240968 473056
rect 235960 473016 235966 473028
rect 240962 473016 240968 473028
rect 241020 473016 241026 473068
rect 216582 472744 216588 472796
rect 216640 472784 216646 472796
rect 235534 472784 235540 472796
rect 216640 472756 235540 472784
rect 216640 472744 216646 472756
rect 235534 472744 235540 472756
rect 235592 472744 235598 472796
rect 32398 472676 32404 472728
rect 32456 472716 32462 472728
rect 224310 472716 224316 472728
rect 32456 472688 224316 472716
rect 32456 472676 32462 472688
rect 224310 472676 224316 472688
rect 224368 472676 224374 472728
rect 235994 472676 236000 472728
rect 236052 472716 236058 472728
rect 324314 472716 324320 472728
rect 236052 472688 324320 472716
rect 236052 472676 236058 472688
rect 324314 472676 324320 472688
rect 324372 472676 324378 472728
rect 215386 472608 215392 472660
rect 215444 472648 215450 472660
rect 511258 472648 511264 472660
rect 215444 472620 511264 472648
rect 215444 472608 215450 472620
rect 511258 472608 511264 472620
rect 511316 472608 511322 472660
rect 40678 471248 40684 471300
rect 40736 471288 40742 471300
rect 224494 471288 224500 471300
rect 40736 471260 224500 471288
rect 40736 471248 40742 471260
rect 224494 471248 224500 471260
rect 224552 471248 224558 471300
rect 237466 471248 237472 471300
rect 237524 471288 237530 471300
rect 440234 471288 440240 471300
rect 237524 471260 440240 471288
rect 237524 471248 237530 471260
rect 440234 471248 440240 471260
rect 440292 471248 440298 471300
rect 214006 470568 214012 470620
rect 214064 470608 214070 470620
rect 579982 470608 579988 470620
rect 214064 470580 579988 470608
rect 214064 470568 214070 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 10318 469888 10324 469940
rect 10376 469928 10382 469940
rect 224678 469928 224684 469940
rect 10376 469900 224684 469928
rect 10376 469888 10382 469900
rect 224678 469888 224684 469900
rect 224736 469888 224742 469940
rect 240318 469888 240324 469940
rect 240376 469928 240382 469940
rect 455414 469928 455420 469940
rect 240376 469900 455420 469928
rect 240376 469888 240382 469900
rect 455414 469888 455420 469900
rect 455472 469888 455478 469940
rect 217318 469820 217324 469872
rect 217376 469860 217382 469872
rect 509878 469860 509884 469872
rect 217376 469832 509884 469860
rect 217376 469820 217382 469832
rect 509878 469820 509884 469832
rect 509936 469820 509942 469872
rect 219618 468596 219624 468648
rect 219676 468636 219682 468648
rect 296070 468636 296076 468648
rect 219676 468608 296076 468636
rect 219676 468596 219682 468608
rect 296070 468596 296076 468608
rect 296128 468596 296134 468648
rect 218330 468528 218336 468580
rect 218388 468568 218394 468580
rect 399478 468568 399484 468580
rect 218388 468540 399484 468568
rect 218388 468528 218394 468540
rect 399478 468528 399484 468540
rect 399536 468528 399542 468580
rect 22738 468460 22744 468512
rect 22796 468500 22802 468512
rect 223758 468500 223764 468512
rect 22796 468472 223764 468500
rect 22796 468460 22802 468472
rect 223758 468460 223764 468472
rect 223816 468460 223822 468512
rect 239030 468460 239036 468512
rect 239088 468500 239094 468512
rect 449894 468500 449900 468512
rect 239088 468472 449900 468500
rect 239088 468460 239094 468472
rect 449894 468460 449900 468472
rect 449952 468460 449958 468512
rect 178678 467236 178684 467288
rect 178736 467276 178742 467288
rect 221366 467276 221372 467288
rect 178736 467248 221372 467276
rect 178736 467236 178742 467248
rect 221366 467236 221372 467248
rect 221424 467236 221430 467288
rect 218422 467168 218428 467220
rect 218480 467208 218486 467220
rect 409138 467208 409144 467220
rect 218480 467180 409144 467208
rect 218480 467168 218486 467180
rect 409138 467168 409144 467180
rect 409196 467168 409202 467220
rect 121362 467100 121368 467152
rect 121420 467140 121426 467152
rect 239490 467140 239496 467152
rect 121420 467112 239496 467140
rect 121420 467100 121426 467112
rect 239490 467100 239496 467112
rect 239548 467100 239554 467152
rect 244550 467100 244556 467152
rect 244608 467140 244614 467152
rect 470594 467140 470600 467152
rect 244608 467112 470600 467140
rect 244608 467100 244614 467112
rect 470594 467100 470600 467112
rect 470652 467100 470658 467152
rect 136542 465808 136548 465860
rect 136600 465848 136606 465860
rect 243354 465848 243360 465860
rect 136600 465820 243360 465848
rect 136600 465808 136606 465820
rect 243354 465808 243360 465820
rect 243412 465808 243418 465860
rect 217502 465740 217508 465792
rect 217560 465780 217566 465792
rect 406378 465780 406384 465792
rect 217560 465752 406384 465780
rect 217560 465740 217566 465752
rect 406378 465740 406384 465752
rect 406436 465740 406442 465792
rect 243078 465672 243084 465724
rect 243136 465712 243142 465724
rect 436738 465712 436744 465724
rect 243136 465684 436744 465712
rect 243136 465672 243142 465684
rect 436738 465672 436744 465684
rect 436796 465672 436802 465724
rect 231486 464448 231492 464500
rect 231544 464488 231550 464500
rect 311894 464488 311900 464500
rect 231544 464460 311900 464488
rect 231544 464448 231550 464460
rect 311894 464448 311900 464460
rect 311952 464448 311958 464500
rect 4062 464380 4068 464432
rect 4120 464420 4126 464432
rect 224218 464420 224224 464432
rect 4120 464392 224224 464420
rect 4120 464380 4126 464392
rect 224218 464380 224224 464392
rect 224276 464380 224282 464432
rect 239214 464380 239220 464432
rect 239272 464420 239278 464432
rect 444374 464420 444380 464432
rect 239272 464392 444380 464420
rect 239272 464380 239278 464392
rect 444374 464380 444380 464392
rect 444432 464380 444438 464432
rect 215846 464312 215852 464364
rect 215904 464352 215910 464364
rect 504358 464352 504364 464364
rect 215904 464324 504364 464352
rect 215904 464312 215910 464324
rect 504358 464312 504364 464324
rect 504416 464312 504422 464364
rect 219710 463156 219716 463208
rect 219768 463196 219774 463208
rect 282914 463196 282920 463208
rect 219768 463168 282920 463196
rect 219768 463156 219774 463168
rect 282914 463156 282920 463168
rect 282972 463156 282978 463208
rect 240502 463088 240508 463140
rect 240560 463128 240566 463140
rect 345014 463128 345020 463140
rect 240560 463100 345020 463128
rect 240560 463088 240566 463100
rect 345014 463088 345020 463100
rect 345072 463088 345078 463140
rect 230750 463020 230756 463072
rect 230808 463060 230814 463072
rect 408034 463060 408040 463072
rect 230808 463032 408040 463060
rect 230808 463020 230814 463032
rect 408034 463020 408040 463032
rect 408092 463020 408098 463072
rect 216858 462952 216864 463004
rect 216916 462992 216922 463004
rect 508498 462992 508504 463004
rect 216916 462964 508504 462992
rect 216916 462952 216922 462964
rect 508498 462952 508504 462964
rect 508556 462952 508562 463004
rect 2866 462340 2872 462392
rect 2924 462380 2930 462392
rect 225598 462380 225604 462392
rect 2924 462352 225604 462380
rect 2924 462340 2930 462352
rect 225598 462340 225604 462352
rect 225656 462340 225662 462392
rect 219894 461796 219900 461848
rect 219952 461836 219958 461848
rect 291838 461836 291844 461848
rect 219952 461808 291844 461836
rect 219952 461796 219958 461808
rect 291838 461796 291844 461808
rect 291896 461796 291902 461848
rect 131022 461728 131028 461780
rect 131080 461768 131086 461780
rect 242066 461768 242072 461780
rect 131080 461740 242072 461768
rect 131080 461728 131086 461740
rect 242066 461728 242072 461740
rect 242124 461728 242130 461780
rect 71774 461660 71780 461712
rect 71832 461700 71838 461712
rect 221550 461700 221556 461712
rect 71832 461672 221556 461700
rect 71832 461660 71838 461672
rect 221550 461660 221556 461672
rect 221608 461660 221614 461712
rect 241790 461660 241796 461712
rect 241848 461700 241854 461712
rect 349154 461700 349160 461712
rect 241848 461672 349160 461700
rect 241848 461660 241854 461672
rect 349154 461660 349160 461672
rect 349212 461660 349218 461712
rect 215754 461592 215760 461644
rect 215812 461632 215818 461644
rect 507118 461632 507124 461644
rect 215812 461604 507124 461632
rect 215812 461592 215818 461604
rect 507118 461592 507124 461604
rect 507176 461592 507182 461644
rect 207658 460844 207664 460896
rect 207716 460884 207722 460896
rect 236546 460884 236552 460896
rect 207716 460856 236552 460884
rect 207716 460844 207722 460856
rect 236546 460844 236552 460856
rect 236604 460844 236610 460896
rect 218606 460300 218612 460352
rect 218664 460340 218670 460352
rect 293218 460340 293224 460352
rect 218664 460312 293224 460340
rect 218664 460300 218670 460312
rect 293218 460300 293224 460312
rect 293276 460300 293282 460352
rect 14458 460232 14464 460284
rect 14516 460272 14522 460284
rect 224034 460272 224040 460284
rect 14516 460244 224040 460272
rect 14516 460232 14522 460244
rect 224034 460232 224040 460244
rect 224092 460232 224098 460284
rect 245838 460232 245844 460284
rect 245896 460272 245902 460284
rect 406470 460272 406476 460284
rect 245896 460244 406476 460272
rect 245896 460232 245902 460244
rect 406470 460232 406476 460244
rect 406528 460232 406534 460284
rect 214190 460164 214196 460216
rect 214248 460204 214254 460216
rect 502978 460204 502984 460216
rect 214248 460176 502984 460204
rect 214248 460164 214254 460176
rect 502978 460164 502984 460176
rect 503036 460164 503042 460216
rect 210418 459484 210424 459536
rect 210476 459524 210482 459536
rect 239122 459524 239128 459536
rect 210476 459496 239128 459524
rect 210476 459484 210482 459496
rect 239122 459484 239128 459496
rect 239180 459524 239186 459536
rect 239398 459524 239404 459536
rect 239180 459496 239404 459524
rect 239180 459484 239186 459496
rect 239398 459484 239404 459496
rect 239456 459484 239462 459536
rect 203518 459416 203524 459468
rect 203576 459456 203582 459468
rect 231578 459456 231584 459468
rect 203576 459428 231584 459456
rect 203576 459416 203582 459428
rect 231578 459416 231584 459428
rect 231636 459416 231642 459468
rect 299658 458940 299664 458992
rect 299716 458980 299722 458992
rect 321278 458980 321284 458992
rect 299716 458952 321284 458980
rect 299716 458940 299722 458952
rect 321278 458940 321284 458952
rect 321336 458940 321342 458992
rect 171962 458872 171968 458924
rect 172020 458912 172026 458924
rect 249794 458912 249800 458924
rect 172020 458884 249800 458912
rect 172020 458872 172026 458884
rect 249794 458872 249800 458884
rect 249852 458872 249858 458924
rect 251818 458872 251824 458924
rect 251876 458912 251882 458924
rect 371510 458912 371516 458924
rect 251876 458884 371516 458912
rect 251876 458872 251882 458884
rect 371510 458872 371516 458884
rect 371568 458872 371574 458924
rect 40034 458804 40040 458856
rect 40092 458844 40098 458856
rect 220998 458844 221004 458856
rect 40092 458816 221004 458844
rect 40092 458804 40098 458816
rect 220998 458804 221004 458816
rect 221056 458804 221062 458856
rect 247034 458804 247040 458856
rect 247092 458844 247098 458856
rect 379882 458844 379888 458856
rect 247092 458816 379888 458844
rect 247092 458804 247098 458816
rect 379882 458804 379888 458816
rect 379940 458804 379946 458856
rect 299382 458736 299388 458788
rect 299440 458776 299446 458788
rect 329650 458776 329656 458788
rect 299440 458748 329656 458776
rect 299440 458736 299446 458748
rect 329650 458736 329656 458748
rect 329708 458736 329714 458788
rect 299474 458668 299480 458720
rect 299532 458708 299538 458720
rect 342530 458708 342536 458720
rect 299532 458680 342536 458708
rect 299532 458668 299538 458680
rect 342530 458668 342536 458680
rect 342588 458668 342594 458720
rect 296070 458600 296076 458652
rect 296128 458640 296134 458652
rect 346394 458640 346400 458652
rect 296128 458612 346400 458640
rect 296128 458600 296134 458612
rect 346394 458600 346400 458612
rect 346452 458600 346458 458652
rect 299566 458532 299572 458584
rect 299624 458572 299630 458584
rect 350902 458572 350908 458584
rect 299624 458544 350908 458572
rect 299624 458532 299630 458544
rect 350902 458532 350908 458544
rect 350960 458532 350966 458584
rect 298922 458464 298928 458516
rect 298980 458504 298986 458516
rect 359274 458504 359280 458516
rect 298980 458476 359280 458504
rect 298980 458464 298986 458476
rect 359274 458464 359280 458476
rect 359332 458464 359338 458516
rect 298002 458396 298008 458448
rect 298060 458436 298066 458448
rect 367646 458436 367652 458448
rect 298060 458408 367652 458436
rect 298060 458396 298066 458408
rect 367646 458396 367652 458408
rect 367704 458396 367710 458448
rect 246298 458328 246304 458380
rect 246356 458368 246362 458380
rect 363138 458368 363144 458380
rect 246356 458340 363144 458368
rect 246356 458328 246362 458340
rect 363138 458328 363144 458340
rect 363196 458328 363202 458380
rect 293310 458260 293316 458312
rect 293368 458300 293374 458312
rect 309042 458300 309048 458312
rect 293368 458272 309048 458300
rect 293368 458260 293374 458272
rect 309042 458260 309048 458272
rect 309100 458260 309106 458312
rect 355962 458192 355968 458244
rect 356020 458232 356026 458244
rect 376018 458232 376024 458244
rect 356020 458204 376024 458232
rect 356020 458192 356026 458204
rect 376018 458192 376024 458204
rect 376076 458192 376082 458244
rect 174538 457512 174544 457564
rect 174596 457552 174602 457564
rect 220814 457552 220820 457564
rect 174596 457524 220820 457552
rect 174596 457512 174602 457524
rect 220814 457512 220820 457524
rect 220872 457512 220878 457564
rect 6914 457444 6920 457496
rect 6972 457484 6978 457496
rect 222010 457484 222016 457496
rect 6972 457456 222016 457484
rect 6972 457444 6978 457456
rect 222010 457444 222016 457456
rect 222068 457444 222074 457496
rect 227346 457444 227352 457496
rect 227404 457484 227410 457496
rect 355962 457484 355968 457496
rect 227404 457456 355968 457484
rect 227404 457444 227410 457456
rect 355962 457444 355968 457456
rect 356020 457444 356026 457496
rect 222930 457240 222936 457292
rect 222988 457280 222994 457292
rect 317414 457280 317420 457292
rect 222988 457252 317420 457280
rect 222988 457240 222994 457252
rect 317414 457240 317420 457252
rect 317472 457240 317478 457292
rect 228450 457172 228456 457224
rect 228508 457212 228514 457224
rect 325786 457212 325792 457224
rect 228508 457184 325792 457212
rect 228508 457172 228514 457184
rect 325786 457172 325792 457184
rect 325844 457172 325850 457224
rect 236362 457104 236368 457156
rect 236420 457144 236426 457156
rect 338022 457144 338028 457156
rect 236420 457116 338028 457144
rect 236420 457104 236426 457116
rect 338022 457104 338028 457116
rect 338080 457104 338086 457156
rect 228542 457036 228548 457088
rect 228600 457076 228606 457088
rect 334158 457076 334164 457088
rect 228600 457048 334164 457076
rect 228600 457036 228606 457048
rect 334158 457036 334164 457048
rect 334216 457036 334222 457088
rect 247126 456968 247132 457020
rect 247184 457008 247190 457020
rect 354766 457008 354772 457020
rect 247184 456980 354772 457008
rect 247184 456968 247190 456980
rect 354766 456968 354772 456980
rect 354824 456968 354830 457020
rect 223022 456900 223028 456952
rect 223080 456940 223086 456952
rect 383746 456940 383752 456952
rect 223080 456912 383752 456940
rect 223080 456900 223086 456912
rect 383746 456900 383752 456912
rect 383804 456900 383810 456952
rect 385310 456872 385316 456884
rect 229066 456844 385316 456872
rect 223850 456764 223856 456816
rect 223908 456804 223914 456816
rect 224310 456804 224316 456816
rect 223908 456776 224316 456804
rect 223908 456764 223914 456776
rect 224310 456764 224316 456776
rect 224368 456804 224374 456816
rect 229066 456804 229094 456844
rect 385310 456832 385316 456844
rect 385368 456832 385374 456884
rect 224368 456776 229094 456804
rect 224368 456764 224374 456776
rect 299014 456764 299020 456816
rect 299072 456804 299078 456816
rect 580166 456804 580172 456816
rect 299072 456776 580172 456804
rect 299072 456764 299078 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 299750 456016 299756 456068
rect 299808 456056 299814 456068
rect 300762 456056 300768 456068
rect 299808 456028 300768 456056
rect 299808 456016 299814 456028
rect 300762 456016 300768 456028
rect 300820 456016 300826 456068
rect 235074 455948 235080 456000
rect 235132 455988 235138 456000
rect 312630 455988 312636 456000
rect 235132 455960 312636 455988
rect 235132 455948 235138 455960
rect 312630 455948 312636 455960
rect 312688 455948 312694 456000
rect 252738 455880 252744 455932
rect 252796 455920 252802 455932
rect 385126 455920 385132 455932
rect 252796 455892 385132 455920
rect 252796 455880 252802 455892
rect 385126 455880 385132 455892
rect 385184 455880 385190 455932
rect 251910 455812 251916 455864
rect 251968 455852 251974 455864
rect 385218 455852 385224 455864
rect 251968 455824 385224 455852
rect 251968 455812 251974 455824
rect 385218 455812 385224 455824
rect 385276 455812 385282 455864
rect 250530 455744 250536 455796
rect 250588 455784 250594 455796
rect 384114 455784 384120 455796
rect 250588 455756 384120 455784
rect 250588 455744 250594 455756
rect 384114 455744 384120 455756
rect 384172 455744 384178 455796
rect 244458 455676 244464 455728
rect 244516 455716 244522 455728
rect 384206 455716 384212 455728
rect 244516 455688 384212 455716
rect 244516 455676 244522 455688
rect 384206 455676 384212 455688
rect 384264 455676 384270 455728
rect 298830 455608 298836 455660
rect 298888 455648 298894 455660
rect 300302 455648 300308 455660
rect 298888 455620 300308 455648
rect 298888 455608 298894 455620
rect 300302 455608 300308 455620
rect 300360 455608 300366 455660
rect 300762 455608 300768 455660
rect 300820 455648 300826 455660
rect 385034 455648 385040 455660
rect 300820 455620 385040 455648
rect 300820 455608 300826 455620
rect 385034 455608 385040 455620
rect 385092 455608 385098 455660
rect 237742 455540 237748 455592
rect 237800 455580 237806 455592
rect 384022 455580 384028 455592
rect 237800 455552 384028 455580
rect 237800 455540 237806 455552
rect 384022 455540 384028 455552
rect 384080 455540 384086 455592
rect 214282 455472 214288 455524
rect 214340 455512 214346 455524
rect 384298 455512 384304 455524
rect 214340 455484 384304 455512
rect 214340 455472 214346 455484
rect 384298 455472 384304 455484
rect 384356 455472 384362 455524
rect 214466 455404 214472 455456
rect 214524 455444 214530 455456
rect 580258 455444 580264 455456
rect 214524 455416 580264 455444
rect 214524 455404 214530 455416
rect 580258 455404 580264 455416
rect 580316 455404 580322 455456
rect 299842 455336 299848 455388
rect 299900 455376 299906 455388
rect 304166 455376 304172 455388
rect 299900 455348 304172 455376
rect 299900 455336 299906 455348
rect 304166 455336 304172 455348
rect 304224 455336 304230 455388
rect 249242 454860 249248 454912
rect 249300 454900 249306 454912
rect 299842 454900 299848 454912
rect 249300 454872 299848 454900
rect 249300 454860 249306 454872
rect 299842 454860 299848 454872
rect 299900 454860 299906 454912
rect 235350 454792 235356 454844
rect 235408 454832 235414 454844
rect 299566 454832 299572 454844
rect 235408 454804 299572 454832
rect 235408 454792 235414 454804
rect 299566 454792 299572 454804
rect 299624 454792 299630 454844
rect 235258 454724 235264 454776
rect 235316 454764 235322 454776
rect 299474 454764 299480 454776
rect 235316 454736 299480 454764
rect 235316 454724 235322 454736
rect 299474 454724 299480 454736
rect 299532 454724 299538 454776
rect 219066 454656 219072 454708
rect 219124 454696 219130 454708
rect 295978 454696 295984 454708
rect 219124 454668 295984 454696
rect 219124 454656 219130 454668
rect 295978 454656 295984 454668
rect 296036 454656 296042 454708
rect 182818 453432 182824 453484
rect 182876 453472 182882 453484
rect 221734 453472 221740 453484
rect 182876 453444 221740 453472
rect 182876 453432 182882 453444
rect 221734 453432 221740 453444
rect 221792 453432 221798 453484
rect 215938 453364 215944 453416
rect 215996 453404 216002 453416
rect 285030 453404 285036 453416
rect 215996 453376 285036 453404
rect 215996 453364 216002 453376
rect 285030 453364 285036 453376
rect 285088 453364 285094 453416
rect 214650 453296 214656 453348
rect 214708 453336 214714 453348
rect 299014 453336 299020 453348
rect 214708 453308 299020 453336
rect 214708 453296 214714 453308
rect 299014 453296 299020 453308
rect 299072 453296 299078 453348
rect 237558 452548 237564 452600
rect 237616 452588 237622 452600
rect 237834 452588 237840 452600
rect 237616 452560 237840 452588
rect 237616 452548 237622 452560
rect 237834 452548 237840 452560
rect 237892 452548 237898 452600
rect 243170 452344 243176 452396
rect 243228 452384 243234 452396
rect 247034 452384 247040 452396
rect 243228 452356 247040 452384
rect 243228 452344 243234 452356
rect 247034 452344 247040 452356
rect 247092 452344 247098 452396
rect 219710 452276 219716 452328
rect 219768 452316 219774 452328
rect 219986 452316 219992 452328
rect 219768 452288 219992 452316
rect 219768 452276 219774 452288
rect 219986 452276 219992 452288
rect 220044 452276 220050 452328
rect 255866 452276 255872 452328
rect 255924 452316 255930 452328
rect 284386 452316 284392 452328
rect 255924 452288 284392 452316
rect 255924 452276 255930 452288
rect 284386 452276 284392 452288
rect 284444 452276 284450 452328
rect 254578 452208 254584 452260
rect 254636 452248 254642 452260
rect 284478 452248 284484 452260
rect 254636 452220 284484 452248
rect 254636 452208 254642 452220
rect 284478 452208 284484 452220
rect 284536 452208 284542 452260
rect 253290 452140 253296 452192
rect 253348 452180 253354 452192
rect 284570 452180 284576 452192
rect 253348 452152 284576 452180
rect 253348 452140 253354 452152
rect 284570 452140 284576 452152
rect 284628 452140 284634 452192
rect 247310 452072 247316 452124
rect 247368 452112 247374 452124
rect 281534 452112 281540 452124
rect 247368 452084 281540 452112
rect 247368 452072 247374 452084
rect 281534 452072 281540 452084
rect 281592 452072 281598 452124
rect 246022 452004 246028 452056
rect 246080 452044 246086 452056
rect 281074 452044 281080 452056
rect 246080 452016 281080 452044
rect 246080 452004 246086 452016
rect 281074 452004 281080 452016
rect 281132 452004 281138 452056
rect 171778 451936 171784 451988
rect 171836 451976 171842 451988
rect 220722 451976 220728 451988
rect 171836 451948 220728 451976
rect 171836 451936 171842 451948
rect 220722 451936 220728 451948
rect 220780 451936 220786 451988
rect 234614 451936 234620 451988
rect 234672 451976 234678 451988
rect 235626 451976 235632 451988
rect 234672 451948 235632 451976
rect 234672 451936 234678 451948
rect 235626 451936 235632 451948
rect 235684 451936 235690 451988
rect 239030 451936 239036 451988
rect 239088 451976 239094 451988
rect 240042 451976 240048 451988
rect 239088 451948 240048 451976
rect 239088 451936 239094 451948
rect 240042 451936 240048 451948
rect 240100 451936 240106 451988
rect 240318 451936 240324 451988
rect 240376 451976 240382 451988
rect 241330 451976 241336 451988
rect 240376 451948 241336 451976
rect 240376 451936 240382 451948
rect 241330 451936 241336 451948
rect 241388 451936 241394 451988
rect 247770 451936 247776 451988
rect 247828 451976 247834 451988
rect 299382 451976 299388 451988
rect 247828 451948 299388 451976
rect 247828 451936 247834 451948
rect 299382 451936 299388 451948
rect 299440 451936 299446 451988
rect 217318 451868 217324 451920
rect 217376 451908 217382 451920
rect 286318 451908 286324 451920
rect 217376 451880 286324 451908
rect 217376 451868 217382 451880
rect 286318 451868 286324 451880
rect 286376 451868 286382 451920
rect 214834 451256 214840 451308
rect 214892 451296 214898 451308
rect 221458 451296 221464 451308
rect 214892 451268 221464 451296
rect 214892 451256 214898 451268
rect 221458 451256 221464 451268
rect 221516 451256 221522 451308
rect 233970 451256 233976 451308
rect 234028 451296 234034 451308
rect 297634 451296 297640 451308
rect 234028 451268 297640 451296
rect 234028 451256 234034 451268
rect 297634 451256 297640 451268
rect 297692 451256 297698 451308
rect 228358 451188 228364 451240
rect 228416 451228 228422 451240
rect 244274 451228 244280 451240
rect 228416 451200 244280 451228
rect 228416 451188 228422 451200
rect 244274 451188 244280 451200
rect 244332 451188 244338 451240
rect 189074 450916 189080 450968
rect 189132 450956 189138 450968
rect 230842 450956 230848 450968
rect 189132 450928 230848 450956
rect 189132 450916 189138 450928
rect 230842 450916 230848 450928
rect 230900 450916 230906 450968
rect 188430 450848 188436 450900
rect 188488 450888 188494 450900
rect 234246 450888 234252 450900
rect 188488 450860 234252 450888
rect 188488 450848 188494 450860
rect 234246 450848 234252 450860
rect 234304 450848 234310 450900
rect 187510 450780 187516 450832
rect 187568 450820 187574 450832
rect 233418 450820 233424 450832
rect 187568 450792 233424 450820
rect 187568 450780 187574 450792
rect 233418 450780 233424 450792
rect 233476 450780 233482 450832
rect 256050 450780 256056 450832
rect 256108 450820 256114 450832
rect 293310 450820 293316 450832
rect 256108 450792 293316 450820
rect 256108 450780 256114 450792
rect 293310 450780 293316 450792
rect 293368 450780 293374 450832
rect 187234 450712 187240 450764
rect 187292 450752 187298 450764
rect 233786 450752 233792 450764
rect 187292 450724 233792 450752
rect 187292 450712 187298 450724
rect 233786 450712 233792 450724
rect 233844 450712 233850 450764
rect 254762 450712 254768 450764
rect 254820 450752 254826 450764
rect 298002 450752 298008 450764
rect 254820 450724 298008 450752
rect 254820 450712 254826 450724
rect 298002 450712 298008 450724
rect 298060 450712 298066 450764
rect 187326 450644 187332 450696
rect 187384 450684 187390 450696
rect 234062 450684 234068 450696
rect 187384 450656 234068 450684
rect 187384 450644 187390 450656
rect 234062 450644 234068 450656
rect 234120 450644 234126 450696
rect 244274 450644 244280 450696
rect 244332 450684 244338 450696
rect 244918 450684 244924 450696
rect 244332 450656 244924 450684
rect 244332 450644 244338 450656
rect 244918 450644 244924 450656
rect 244976 450644 244982 450696
rect 255682 450644 255688 450696
rect 255740 450684 255746 450696
rect 299750 450684 299756 450696
rect 255740 450656 299756 450684
rect 255740 450644 255746 450656
rect 299750 450644 299756 450656
rect 299808 450644 299814 450696
rect 187418 450576 187424 450628
rect 187476 450616 187482 450628
rect 255406 450616 255412 450628
rect 187476 450588 255412 450616
rect 187476 450576 187482 450588
rect 255406 450576 255412 450588
rect 255464 450576 255470 450628
rect 187602 450508 187608 450560
rect 187660 450548 187666 450560
rect 255314 450548 255320 450560
rect 187660 450520 255320 450548
rect 187660 450508 187666 450520
rect 255314 450508 255320 450520
rect 255372 450508 255378 450560
rect 230106 449896 230112 449948
rect 230164 449936 230170 449948
rect 293218 449936 293224 449948
rect 230164 449908 293224 449936
rect 230164 449896 230170 449908
rect 293218 449896 293224 449908
rect 293276 449896 293282 449948
rect 3510 449828 3516 449880
rect 3568 449868 3574 449880
rect 223022 449868 223028 449880
rect 3568 449840 223028 449868
rect 3568 449828 3574 449840
rect 223022 449828 223028 449840
rect 223080 449828 223086 449880
rect 234246 449828 234252 449880
rect 234304 449868 234310 449880
rect 234522 449868 234528 449880
rect 234304 449840 234528 449868
rect 234304 449828 234310 449840
rect 234522 449828 234528 449840
rect 234580 449868 234586 449880
rect 297174 449868 297180 449880
rect 234580 449840 297180 449868
rect 234580 449828 234586 449840
rect 297174 449828 297180 449840
rect 297232 449828 297238 449880
rect 229738 449760 229744 449812
rect 229796 449800 229802 449812
rect 242986 449800 242992 449812
rect 229796 449772 242992 449800
rect 229796 449760 229802 449772
rect 242986 449760 242992 449772
rect 243044 449800 243050 449812
rect 243538 449800 243544 449812
rect 243044 449772 243544 449800
rect 243044 449760 243050 449772
rect 243538 449760 243544 449772
rect 243596 449760 243602 449812
rect 253842 449760 253848 449812
rect 253900 449800 253906 449812
rect 281810 449800 281816 449812
rect 253900 449772 281816 449800
rect 253900 449760 253906 449772
rect 281810 449760 281816 449772
rect 281868 449760 281874 449812
rect 187142 449692 187148 449744
rect 187200 449732 187206 449744
rect 232682 449732 232688 449744
rect 187200 449704 232688 449732
rect 187200 449692 187206 449704
rect 232682 449692 232688 449704
rect 232740 449692 232746 449744
rect 252554 449692 252560 449744
rect 252612 449732 252618 449744
rect 282086 449732 282092 449744
rect 252612 449704 282092 449732
rect 252612 449692 252618 449704
rect 282086 449692 282092 449704
rect 282144 449692 282150 449744
rect 189902 449624 189908 449676
rect 189960 449664 189966 449676
rect 247402 449664 247408 449676
rect 189960 449636 247408 449664
rect 189960 449624 189966 449636
rect 247402 449624 247408 449636
rect 247460 449624 247466 449676
rect 251266 449624 251272 449676
rect 251324 449664 251330 449676
rect 281902 449664 281908 449676
rect 251324 449636 281908 449664
rect 251324 449624 251330 449636
rect 281902 449624 281908 449636
rect 281960 449624 281966 449676
rect 189994 449556 190000 449608
rect 190052 449596 190058 449608
rect 246114 449596 246120 449608
rect 190052 449568 246120 449596
rect 190052 449556 190058 449568
rect 246114 449556 246120 449568
rect 246172 449556 246178 449608
rect 249978 449556 249984 449608
rect 250036 449596 250042 449608
rect 281994 449596 282000 449608
rect 250036 449568 282000 449596
rect 250036 449556 250042 449568
rect 281994 449556 282000 449568
rect 282052 449556 282058 449608
rect 188338 449488 188344 449540
rect 188396 449528 188402 449540
rect 247218 449528 247224 449540
rect 188396 449500 247224 449528
rect 188396 449488 188402 449500
rect 247218 449488 247224 449500
rect 247276 449488 247282 449540
rect 250714 449488 250720 449540
rect 250772 449528 250778 449540
rect 283190 449528 283196 449540
rect 250772 449500 283196 449528
rect 250772 449488 250778 449500
rect 283190 449488 283196 449500
rect 283248 449488 283254 449540
rect 252002 449420 252008 449472
rect 252060 449460 252066 449472
rect 284294 449460 284300 449472
rect 252060 449432 284300 449460
rect 252060 449420 252066 449432
rect 284294 449420 284300 449432
rect 284352 449420 284358 449472
rect 140682 449352 140688 449404
rect 140740 449392 140746 449404
rect 244642 449392 244648 449404
rect 140740 449364 244648 449392
rect 140740 449352 140746 449364
rect 244642 449352 244648 449364
rect 244700 449352 244706 449404
rect 248690 449352 248696 449404
rect 248748 449392 248754 449404
rect 281626 449392 281632 449404
rect 248748 449364 281632 449392
rect 248748 449352 248754 449364
rect 281626 449352 281632 449364
rect 281684 449352 281690 449404
rect 115842 449284 115848 449336
rect 115900 449324 115906 449336
rect 238202 449324 238208 449336
rect 115900 449296 238208 449324
rect 115900 449284 115906 449296
rect 238202 449284 238208 449296
rect 238260 449284 238266 449336
rect 249426 449284 249432 449336
rect 249484 449324 249490 449336
rect 283098 449324 283104 449336
rect 249484 449296 283104 449324
rect 249484 449284 249490 449296
rect 283098 449284 283104 449296
rect 283156 449284 283162 449336
rect 111702 449216 111708 449268
rect 111760 449256 111766 449268
rect 236914 449256 236920 449268
rect 111760 449228 236920 449256
rect 111760 449216 111766 449228
rect 236914 449216 236920 449228
rect 236972 449216 236978 449268
rect 246758 449216 246764 449268
rect 246816 449256 246822 449268
rect 298922 449256 298928 449268
rect 246816 449228 298928 449256
rect 246816 449216 246822 449228
rect 298922 449216 298928 449228
rect 298980 449216 298986 449268
rect 3878 449148 3884 449200
rect 3936 449188 3942 449200
rect 223114 449188 223120 449200
rect 3936 449160 223120 449188
rect 3936 449148 3942 449160
rect 223114 449148 223120 449160
rect 223172 449148 223178 449200
rect 241514 449148 241520 449200
rect 241572 449188 241578 449200
rect 298830 449188 298836 449200
rect 241572 449160 298836 449188
rect 241572 449148 241578 449160
rect 298830 449148 298836 449160
rect 298888 449148 298894 449200
rect 204898 449080 204904 449132
rect 204956 449120 204962 449132
rect 232590 449120 232596 449132
rect 204956 449092 232596 449120
rect 204956 449080 204962 449092
rect 232590 449080 232596 449092
rect 232648 449080 232654 449132
rect 255130 449080 255136 449132
rect 255188 449120 255194 449132
rect 281718 449120 281724 449132
rect 255188 449092 281724 449120
rect 255188 449080 255194 449092
rect 281718 449080 281724 449092
rect 281776 449080 281782 449132
rect 186958 449012 186964 449064
rect 187016 449052 187022 449064
rect 233050 449052 233056 449064
rect 187016 449024 233056 449052
rect 187016 449012 187022 449024
rect 233050 449012 233056 449024
rect 233108 449012 233114 449064
rect 171870 448944 171876 448996
rect 171928 448984 171934 448996
rect 252370 448984 252376 448996
rect 171928 448956 252376 448984
rect 171928 448944 171934 448956
rect 252370 448944 252376 448956
rect 252428 448944 252434 448996
rect 252186 448604 252192 448656
rect 252244 448644 252250 448656
rect 293310 448644 293316 448656
rect 252244 448616 293316 448644
rect 252244 448604 252250 448616
rect 293310 448604 293316 448616
rect 293368 448604 293374 448656
rect 222746 448536 222752 448588
rect 222804 448576 222810 448588
rect 223022 448576 223028 448588
rect 222804 448548 223028 448576
rect 222804 448536 222810 448548
rect 223022 448536 223028 448548
rect 223080 448536 223086 448588
rect 247034 448536 247040 448588
rect 247092 448576 247098 448588
rect 293402 448576 293408 448588
rect 247092 448548 293408 448576
rect 247092 448536 247098 448548
rect 293402 448536 293408 448548
rect 293460 448536 293466 448588
rect 23474 448468 23480 448520
rect 23532 448508 23538 448520
rect 222194 448508 222200 448520
rect 23532 448480 222200 448508
rect 23532 448468 23538 448480
rect 222194 448468 222200 448480
rect 222252 448508 222258 448520
rect 222930 448508 222936 448520
rect 222252 448480 222936 448508
rect 222252 448468 222258 448480
rect 222930 448468 222936 448480
rect 222988 448468 222994 448520
rect 297726 448508 297732 448520
rect 234586 448480 297732 448508
rect 233050 448400 233056 448452
rect 233108 448440 233114 448452
rect 234586 448440 234614 448480
rect 297726 448468 297732 448480
rect 297784 448468 297790 448520
rect 297358 448440 297364 448452
rect 233108 448412 234614 448440
rect 239416 448412 297364 448440
rect 233108 448400 233114 448412
rect 222838 448332 222844 448384
rect 222896 448372 222902 448384
rect 231946 448372 231952 448384
rect 222896 448344 231952 448372
rect 222896 448332 222902 448344
rect 231946 448332 231952 448344
rect 232004 448372 232010 448384
rect 232498 448372 232504 448384
rect 232004 448344 232504 448372
rect 232004 448332 232010 448344
rect 232498 448332 232504 448344
rect 232556 448332 232562 448384
rect 232682 448332 232688 448384
rect 232740 448372 232746 448384
rect 239416 448372 239444 448412
rect 297358 448400 297364 448412
rect 297416 448400 297422 448452
rect 232740 448344 239444 448372
rect 232740 448332 232746 448344
rect 240410 448332 240416 448384
rect 240468 448372 240474 448384
rect 240778 448372 240784 448384
rect 240468 448344 240784 448372
rect 240468 448332 240474 448344
rect 240778 448332 240784 448344
rect 240836 448332 240842 448384
rect 297818 448372 297824 448384
rect 240980 448344 297824 448372
rect 233786 448264 233792 448316
rect 233844 448304 233850 448316
rect 239398 448304 239404 448316
rect 233844 448276 239404 448304
rect 233844 448264 233850 448276
rect 239398 448264 239404 448276
rect 239456 448264 239462 448316
rect 184198 448196 184204 448248
rect 184256 448236 184262 448248
rect 221642 448236 221648 448248
rect 184256 448208 221648 448236
rect 184256 448196 184262 448208
rect 221642 448196 221648 448208
rect 221700 448196 221706 448248
rect 226978 448196 226984 448248
rect 227036 448236 227042 448248
rect 240410 448236 240416 448248
rect 227036 448208 240416 448236
rect 227036 448196 227042 448208
rect 240410 448196 240416 448208
rect 240468 448196 240474 448248
rect 3694 448128 3700 448180
rect 3752 448168 3758 448180
rect 222930 448168 222936 448180
rect 3752 448140 222936 448168
rect 3752 448128 3758 448140
rect 222930 448128 222936 448140
rect 222988 448128 222994 448180
rect 233418 448128 233424 448180
rect 233476 448168 233482 448180
rect 240980 448168 241008 448344
rect 297818 448332 297824 448344
rect 297876 448332 297882 448384
rect 297450 448304 297456 448316
rect 248386 448276 297456 448304
rect 248386 448236 248414 448276
rect 297450 448264 297456 448276
rect 297508 448264 297514 448316
rect 233476 448140 241008 448168
rect 244246 448208 248414 448236
rect 233476 448128 233482 448140
rect 3970 448060 3976 448112
rect 4028 448100 4034 448112
rect 223482 448100 223488 448112
rect 4028 448072 223488 448100
rect 4028 448060 4034 448072
rect 223482 448060 223488 448072
rect 223540 448060 223546 448112
rect 239398 448060 239404 448112
rect 239456 448100 239462 448112
rect 244246 448100 244274 448208
rect 255314 448196 255320 448248
rect 255372 448236 255378 448248
rect 256234 448236 256240 448248
rect 255372 448208 256240 448236
rect 255372 448196 255378 448208
rect 256234 448196 256240 448208
rect 256292 448236 256298 448248
rect 297542 448236 297548 448248
rect 256292 448208 297548 448236
rect 256292 448196 256298 448208
rect 297542 448196 297548 448208
rect 297600 448196 297606 448248
rect 239456 448072 244274 448100
rect 239456 448060 239462 448072
rect 3418 447992 3424 448044
rect 3476 448032 3482 448044
rect 222378 448032 222384 448044
rect 3476 448004 222384 448032
rect 3476 447992 3482 448004
rect 222378 447992 222384 448004
rect 222436 447992 222442 448044
rect 3602 447924 3608 447976
rect 3660 447964 3666 447976
rect 222562 447964 222568 447976
rect 3660 447936 222568 447964
rect 3660 447924 3666 447936
rect 222562 447924 222568 447936
rect 222620 447924 222626 447976
rect 236730 447924 236736 447976
rect 236788 447964 236794 447976
rect 251818 447964 251824 447976
rect 236788 447936 251824 447964
rect 236788 447924 236794 447936
rect 251818 447924 251824 447936
rect 251876 447924 251882 447976
rect 3786 447856 3792 447908
rect 3844 447896 3850 447908
rect 223298 447896 223304 447908
rect 3844 447868 223304 447896
rect 3844 447856 3850 447868
rect 223298 447856 223304 447868
rect 223356 447856 223362 447908
rect 231762 447856 231768 447908
rect 231820 447896 231826 447908
rect 239674 447896 239680 447908
rect 231820 447868 239680 447896
rect 231820 447856 231826 447868
rect 239674 447856 239680 447868
rect 239732 447856 239738 447908
rect 248874 447856 248880 447908
rect 248932 447896 248938 447908
rect 280982 447896 280988 447908
rect 248932 447868 280988 447896
rect 248932 447856 248938 447868
rect 280982 447856 280988 447868
rect 281040 447856 281046 447908
rect 3234 447788 3240 447840
rect 3292 447828 3298 447840
rect 224770 447828 224776 447840
rect 3292 447800 224776 447828
rect 3292 447788 3298 447800
rect 224770 447788 224776 447800
rect 224828 447788 224834 447840
rect 226242 447788 226248 447840
rect 226300 447828 226306 447840
rect 238386 447828 238392 447840
rect 226300 447800 238392 447828
rect 226300 447788 226306 447800
rect 238386 447788 238392 447800
rect 238444 447788 238450 447840
rect 245654 447788 245660 447840
rect 245712 447828 245718 447840
rect 296070 447828 296076 447840
rect 245712 447800 296076 447828
rect 245712 447788 245718 447800
rect 296070 447788 296076 447800
rect 296128 447788 296134 447840
rect 213178 447720 213184 447772
rect 213236 447760 213242 447772
rect 219158 447760 219164 447772
rect 213236 447732 219164 447760
rect 213236 447720 213242 447732
rect 219158 447720 219164 447732
rect 219216 447720 219222 447772
rect 245838 447720 245844 447772
rect 245896 447760 245902 447772
rect 246390 447760 246396 447772
rect 245896 447732 246396 447760
rect 245896 447720 245902 447732
rect 246390 447720 246396 447732
rect 246448 447720 246454 447772
rect 211706 447652 211712 447704
rect 211764 447692 211770 447704
rect 218790 447692 218796 447704
rect 211764 447664 218796 447692
rect 211764 447652 211770 447664
rect 218790 447652 218796 447664
rect 218848 447652 218854 447704
rect 219434 447652 219440 447704
rect 219492 447692 219498 447704
rect 219894 447692 219900 447704
rect 219492 447664 219900 447692
rect 219492 447652 219498 447664
rect 219894 447652 219900 447664
rect 219952 447652 219958 447704
rect 246022 447652 246028 447704
rect 246080 447692 246086 447704
rect 246850 447692 246856 447704
rect 246080 447664 246856 447692
rect 246080 447652 246086 447664
rect 246850 447652 246856 447664
rect 246908 447652 246914 447704
rect 212810 447584 212816 447636
rect 212868 447624 212874 447636
rect 212868 447596 219434 447624
rect 212868 447584 212874 447596
rect 212626 447516 212632 447568
rect 212684 447556 212690 447568
rect 212684 447528 219020 447556
rect 212684 447516 212690 447528
rect 212258 447448 212264 447500
rect 212316 447488 212322 447500
rect 212316 447460 216628 447488
rect 212316 447448 212322 447460
rect 214006 447312 214012 447364
rect 214064 447352 214070 447364
rect 215018 447352 215024 447364
rect 214064 447324 215024 447352
rect 214064 447312 214070 447324
rect 215018 447312 215024 447324
rect 215076 447312 215082 447364
rect 215662 447312 215668 447364
rect 215720 447352 215726 447364
rect 216490 447352 216496 447364
rect 215720 447324 216496 447352
rect 215720 447312 215726 447324
rect 216490 447312 216496 447324
rect 216548 447312 216554 447364
rect 214190 447244 214196 447296
rect 214248 447284 214254 447296
rect 215202 447284 215208 447296
rect 214248 447256 215208 447284
rect 214248 447244 214254 447256
rect 215202 447244 215208 447256
rect 215260 447244 215266 447296
rect 215846 447244 215852 447296
rect 215904 447284 215910 447296
rect 216306 447284 216312 447296
rect 215904 447256 216312 447284
rect 215904 447244 215910 447256
rect 216306 447244 216312 447256
rect 216364 447244 216370 447296
rect 215294 447176 215300 447228
rect 215352 447216 215358 447228
rect 216122 447216 216128 447228
rect 215352 447188 216128 447216
rect 215352 447176 215358 447188
rect 216122 447176 216128 447188
rect 216180 447176 216186 447228
rect 216600 447216 216628 447460
rect 217134 447312 217140 447364
rect 217192 447352 217198 447364
rect 217594 447352 217600 447364
rect 217192 447324 217600 447352
rect 217192 447312 217198 447324
rect 217594 447312 217600 447324
rect 217652 447312 217658 447364
rect 218054 447312 218060 447364
rect 218112 447352 218118 447364
rect 218882 447352 218888 447364
rect 218112 447324 218888 447352
rect 218112 447312 218118 447324
rect 218882 447312 218888 447324
rect 218940 447312 218946 447364
rect 218992 447352 219020 447528
rect 219406 447488 219434 447596
rect 241882 447584 241888 447636
rect 241940 447624 241946 447636
rect 246298 447624 246304 447636
rect 241940 447596 246304 447624
rect 241940 447584 241946 447596
rect 246298 447584 246304 447596
rect 246356 447584 246362 447636
rect 220998 447516 221004 447568
rect 221056 447556 221062 447568
rect 221826 447556 221832 447568
rect 221056 447528 221832 447556
rect 221056 447516 221062 447528
rect 221826 447516 221832 447528
rect 221884 447516 221890 447568
rect 240594 447516 240600 447568
rect 240652 447556 240658 447568
rect 298002 447556 298008 447568
rect 240652 447528 298008 447556
rect 240652 447516 240658 447528
rect 298002 447516 298008 447528
rect 298060 447516 298066 447568
rect 296346 447488 296352 447500
rect 219406 447460 296352 447488
rect 296346 447448 296352 447460
rect 296404 447448 296410 447500
rect 219158 447380 219164 447432
rect 219216 447420 219222 447432
rect 296622 447420 296628 447432
rect 219216 447392 296628 447420
rect 219216 447380 219222 447392
rect 296622 447380 296628 447392
rect 296680 447380 296686 447432
rect 296438 447352 296444 447364
rect 218992 447324 296444 447352
rect 296438 447312 296444 447324
rect 296496 447312 296502 447364
rect 218238 447244 218244 447296
rect 218296 447284 218302 447296
rect 218698 447284 218704 447296
rect 218296 447256 218704 447284
rect 218296 447244 218302 447256
rect 218698 447244 218704 447256
rect 218756 447244 218762 447296
rect 218790 447244 218796 447296
rect 218848 447284 218854 447296
rect 296162 447284 296168 447296
rect 218848 447256 296168 447284
rect 218848 447244 218854 447256
rect 296162 447244 296168 447256
rect 296220 447244 296226 447296
rect 296254 447216 296260 447228
rect 216600 447188 296260 447216
rect 296254 447176 296260 447188
rect 296312 447176 296318 447228
rect 213730 447108 213736 447160
rect 213788 447148 213794 447160
rect 299198 447148 299204 447160
rect 213788 447120 299204 447148
rect 213788 447108 213794 447120
rect 299198 447108 299204 447120
rect 299256 447108 299262 447160
rect 232038 447040 232044 447092
rect 232096 447080 232102 447092
rect 232498 447080 232504 447092
rect 232096 447052 232504 447080
rect 232096 447040 232102 447052
rect 232498 447040 232504 447052
rect 232556 447040 232562 447092
rect 252922 447040 252928 447092
rect 252980 447080 252986 447092
rect 282362 447080 282368 447092
rect 252980 447052 282368 447080
rect 252980 447040 252986 447052
rect 282362 447040 282368 447052
rect 282420 447040 282426 447092
rect 255314 446972 255320 447024
rect 255372 447012 255378 447024
rect 286410 447012 286416 447024
rect 255372 446984 286416 447012
rect 255372 446972 255378 446984
rect 286410 446972 286416 446984
rect 286468 446972 286474 447024
rect 250346 446904 250352 446956
rect 250404 446944 250410 446956
rect 282270 446944 282276 446956
rect 250404 446916 282276 446944
rect 250404 446904 250410 446916
rect 282270 446904 282276 446916
rect 282328 446904 282334 446956
rect 224954 446836 224960 446888
rect 225012 446876 225018 446888
rect 225598 446876 225604 446888
rect 225012 446848 225604 446876
rect 225012 446836 225018 446848
rect 225598 446836 225604 446848
rect 225656 446836 225662 446888
rect 243722 446836 243728 446888
rect 243780 446876 243786 446888
rect 246666 446876 246672 446888
rect 243780 446848 246672 446876
rect 243780 446836 243786 446848
rect 246666 446836 246672 446848
rect 246724 446836 246730 446888
rect 247770 446836 247776 446888
rect 247828 446876 247834 446888
rect 282178 446876 282184 446888
rect 247828 446848 282184 446876
rect 247828 446836 247834 446848
rect 282178 446836 282184 446848
rect 282236 446836 282242 446888
rect 3694 446768 3700 446820
rect 3752 446808 3758 446820
rect 227530 446808 227536 446820
rect 3752 446780 227536 446808
rect 3752 446768 3758 446780
rect 227530 446768 227536 446780
rect 227588 446768 227594 446820
rect 250162 446768 250168 446820
rect 250220 446808 250226 446820
rect 284938 446808 284944 446820
rect 250220 446780 284944 446808
rect 250220 446768 250226 446780
rect 284938 446768 284944 446780
rect 284996 446768 285002 446820
rect 221642 446700 221648 446752
rect 221700 446740 221706 446752
rect 248598 446740 248604 446752
rect 221700 446712 248604 446740
rect 221700 446700 221706 446712
rect 248598 446700 248604 446712
rect 248656 446700 248662 446752
rect 251450 446700 251456 446752
rect 251508 446740 251514 446752
rect 289170 446740 289176 446752
rect 251508 446712 289176 446740
rect 251508 446700 251514 446712
rect 289170 446700 289176 446712
rect 289228 446700 289234 446752
rect 3418 446632 3424 446684
rect 3476 446672 3482 446684
rect 228634 446672 228640 446684
rect 3476 446644 228640 446672
rect 3476 446632 3482 446644
rect 228634 446632 228640 446644
rect 228692 446632 228698 446684
rect 252738 446632 252744 446684
rect 252796 446672 252802 446684
rect 291930 446672 291936 446684
rect 252796 446644 291936 446672
rect 252796 446632 252802 446644
rect 291930 446632 291936 446644
rect 291988 446632 291994 446684
rect 4982 446564 4988 446616
rect 5040 446604 5046 446616
rect 225506 446604 225512 446616
rect 5040 446576 225512 446604
rect 5040 446564 5046 446576
rect 225506 446564 225512 446576
rect 225564 446564 225570 446616
rect 246298 446564 246304 446616
rect 246356 446604 246362 446616
rect 287698 446604 287704 446616
rect 246356 446576 287704 446604
rect 246356 446564 246362 446576
rect 287698 446564 287704 446576
rect 287756 446564 287762 446616
rect 216582 446496 216588 446548
rect 216640 446536 216646 446548
rect 227162 446536 227168 446548
rect 216640 446508 227168 446536
rect 216640 446496 216646 446508
rect 227162 446496 227168 446508
rect 227220 446496 227226 446548
rect 247586 446496 247592 446548
rect 247644 446536 247650 446548
rect 289078 446536 289084 446548
rect 247644 446508 289084 446536
rect 247644 446496 247650 446508
rect 289078 446496 289084 446508
rect 289136 446496 289142 446548
rect 188890 446428 188896 446480
rect 188948 446468 188954 446480
rect 220354 446468 220360 446480
rect 188948 446440 220360 446468
rect 188948 446428 188954 446440
rect 220354 446428 220360 446440
rect 220412 446428 220418 446480
rect 238938 446428 238944 446480
rect 238996 446468 239002 446480
rect 243630 446468 243636 446480
rect 238996 446440 243636 446468
rect 238996 446428 239002 446440
rect 243630 446428 243636 446440
rect 243688 446428 243694 446480
rect 244826 446428 244832 446480
rect 244884 446468 244890 446480
rect 252646 446468 252652 446480
rect 244884 446440 252652 446468
rect 244884 446428 244890 446440
rect 252646 446428 252652 446440
rect 252704 446428 252710 446480
rect 256602 446428 256608 446480
rect 256660 446468 256666 446480
rect 299842 446468 299848 446480
rect 256660 446440 299848 446468
rect 256660 446428 256666 446440
rect 299842 446428 299848 446440
rect 299900 446428 299906 446480
rect 188982 446360 188988 446412
rect 189040 446400 189046 446412
rect 220538 446400 220544 446412
rect 189040 446372 220544 446400
rect 189040 446360 189046 446372
rect 220538 446360 220544 446372
rect 220596 446360 220602 446412
rect 229922 446360 229928 446412
rect 229980 446400 229986 446412
rect 230658 446400 230664 446412
rect 229980 446372 230664 446400
rect 229980 446360 229986 446372
rect 230658 446360 230664 446372
rect 230716 446360 230722 446412
rect 233234 446360 233240 446412
rect 233292 446400 233298 446412
rect 251910 446400 251916 446412
rect 233292 446372 251916 446400
rect 233292 446360 233298 446372
rect 251910 446360 251916 446372
rect 251968 446360 251974 446412
rect 254026 446360 254032 446412
rect 254084 446400 254090 446412
rect 298738 446400 298744 446412
rect 254084 446372 298744 446400
rect 254084 446360 254090 446372
rect 298738 446360 298744 446372
rect 298796 446360 298802 446412
rect 212074 446292 212080 446344
rect 212132 446332 212138 446344
rect 299014 446332 299020 446344
rect 212132 446304 299020 446332
rect 212132 446292 212138 446304
rect 299014 446292 299020 446304
rect 299072 446292 299078 446344
rect 213362 446224 213368 446276
rect 213420 446264 213426 446276
rect 296530 446264 296536 446276
rect 213420 446236 296536 446264
rect 213420 446224 213426 446236
rect 296530 446224 296536 446236
rect 296588 446224 296594 446276
rect 214098 446156 214104 446208
rect 214156 446196 214162 446208
rect 298554 446196 298560 446208
rect 214156 446168 298560 446196
rect 214156 446156 214162 446168
rect 298554 446156 298560 446168
rect 298612 446156 298618 446208
rect 4890 446088 4896 446140
rect 4948 446128 4954 446140
rect 226058 446128 226064 446140
rect 4948 446100 226064 446128
rect 4948 446088 4954 446100
rect 226058 446088 226064 446100
rect 226116 446088 226122 446140
rect 234338 446088 234344 446140
rect 234396 446128 234402 446140
rect 255590 446128 255596 446140
rect 234396 446100 255596 446128
rect 234396 446088 234402 446100
rect 255590 446088 255596 446100
rect 255648 446088 255654 446140
rect 3878 446020 3884 446072
rect 3936 446060 3942 446072
rect 226978 446060 226984 446072
rect 3936 446032 226984 446060
rect 3936 446020 3942 446032
rect 226978 446020 226984 446032
rect 227036 446020 227042 446072
rect 231394 446020 231400 446072
rect 231452 446060 231458 446072
rect 255406 446060 255412 446072
rect 231452 446032 255412 446060
rect 231452 446020 231458 446032
rect 255406 446020 255412 446032
rect 255464 446020 255470 446072
rect 224954 445952 224960 446004
rect 225012 445992 225018 446004
rect 254302 445992 254308 446004
rect 225012 445964 254308 445992
rect 225012 445952 225018 445964
rect 254302 445952 254308 445964
rect 254360 445952 254366 446004
rect 4798 445884 4804 445936
rect 4856 445924 4862 445936
rect 228818 445924 228824 445936
rect 4856 445896 228824 445924
rect 4856 445884 4862 445896
rect 228818 445884 228824 445896
rect 228876 445884 228882 445936
rect 239306 445884 239312 445936
rect 239364 445924 239370 445936
rect 239364 445896 243584 445924
rect 239364 445884 239370 445896
rect 3786 445816 3792 445868
rect 3844 445856 3850 445868
rect 227714 445856 227720 445868
rect 3844 445828 227720 445856
rect 3844 445816 3850 445828
rect 227714 445816 227720 445828
rect 227772 445816 227778 445868
rect 229830 445816 229836 445868
rect 229888 445856 229894 445868
rect 237098 445856 237104 445868
rect 229888 445828 237104 445856
rect 229888 445816 229894 445828
rect 237098 445816 237104 445828
rect 237156 445816 237162 445868
rect 242618 445816 242624 445868
rect 242676 445856 242682 445868
rect 243446 445856 243452 445868
rect 242676 445828 243452 445856
rect 242676 445816 242682 445828
rect 243446 445816 243452 445828
rect 243504 445816 243510 445868
rect 243556 445856 243584 445896
rect 243630 445884 243636 445936
rect 243688 445924 243694 445936
rect 244826 445924 244832 445936
rect 243688 445896 244832 445924
rect 243688 445884 243694 445896
rect 244826 445884 244832 445896
rect 244884 445884 244890 445936
rect 249886 445924 249892 445936
rect 244936 445896 249892 445924
rect 244936 445856 244964 445896
rect 249886 445884 249892 445896
rect 249944 445884 249950 445936
rect 243556 445828 244964 445856
rect 245010 445816 245016 445868
rect 245068 445856 245074 445868
rect 248046 445856 248052 445868
rect 245068 445828 248052 445856
rect 245068 445816 245074 445828
rect 248046 445816 248052 445828
rect 248104 445816 248110 445868
rect 219342 445748 219348 445800
rect 219400 445788 219406 445800
rect 225138 445788 225144 445800
rect 219400 445760 225144 445788
rect 219400 445748 219406 445760
rect 225138 445748 225144 445760
rect 225196 445748 225202 445800
rect 232866 445748 232872 445800
rect 232924 445788 232930 445800
rect 232924 445760 244780 445788
rect 232924 445748 232930 445760
rect 227898 445680 227904 445732
rect 227956 445720 227962 445732
rect 228450 445720 228456 445732
rect 227956 445692 228456 445720
rect 227956 445680 227962 445692
rect 228450 445680 228456 445692
rect 228508 445680 228514 445732
rect 244752 445720 244780 445760
rect 244826 445748 244832 445800
rect 244884 445788 244890 445800
rect 246574 445788 246580 445800
rect 244884 445760 246580 445788
rect 244884 445748 244890 445760
rect 246574 445748 246580 445760
rect 246632 445748 246638 445800
rect 245654 445720 245660 445732
rect 244752 445692 245660 445720
rect 245654 445680 245660 445692
rect 245712 445680 245718 445732
rect 211522 445340 211528 445392
rect 211580 445380 211586 445392
rect 220078 445380 220084 445392
rect 211580 445352 220084 445380
rect 211580 445340 211586 445352
rect 220078 445340 220084 445352
rect 220136 445340 220142 445392
rect 221090 445340 221096 445392
rect 221148 445380 221154 445392
rect 221734 445380 221740 445392
rect 221148 445352 221740 445380
rect 221148 445340 221154 445352
rect 221734 445340 221740 445352
rect 221792 445340 221798 445392
rect 247126 445340 247132 445392
rect 247184 445380 247190 445392
rect 248322 445380 248328 445392
rect 247184 445352 248328 445380
rect 247184 445340 247190 445352
rect 248322 445340 248328 445352
rect 248380 445340 248386 445392
rect 196710 445272 196716 445324
rect 196768 445312 196774 445324
rect 226794 445312 226800 445324
rect 196768 445284 226800 445312
rect 196768 445272 196774 445284
rect 226794 445272 226800 445284
rect 226852 445312 226858 445324
rect 226852 445284 229094 445312
rect 226852 445272 226858 445284
rect 98638 445204 98644 445256
rect 98696 445244 98702 445256
rect 225690 445244 225696 445256
rect 98696 445216 225696 445244
rect 98696 445204 98702 445216
rect 225690 445204 225696 445216
rect 225748 445204 225754 445256
rect 229066 445244 229094 445284
rect 229554 445272 229560 445324
rect 229612 445312 229618 445324
rect 266998 445312 267004 445324
rect 229612 445284 267004 445312
rect 229612 445272 229618 445284
rect 266998 445272 267004 445284
rect 267056 445272 267062 445324
rect 265894 445244 265900 445256
rect 229066 445216 265900 445244
rect 265894 445204 265900 445216
rect 265952 445204 265958 445256
rect 199562 445136 199568 445188
rect 199620 445176 199626 445188
rect 226242 445176 226248 445188
rect 199620 445148 226248 445176
rect 199620 445136 199626 445148
rect 226242 445136 226248 445148
rect 226300 445136 226306 445188
rect 234706 445136 234712 445188
rect 234764 445176 234770 445188
rect 235350 445176 235356 445188
rect 234764 445148 235356 445176
rect 234764 445136 234770 445148
rect 235350 445136 235356 445148
rect 235408 445136 235414 445188
rect 236270 445136 236276 445188
rect 236328 445176 236334 445188
rect 237282 445176 237288 445188
rect 236328 445148 237288 445176
rect 236328 445136 236334 445148
rect 237282 445136 237288 445148
rect 237340 445136 237346 445188
rect 238754 445136 238760 445188
rect 238812 445176 238818 445188
rect 239214 445176 239220 445188
rect 238812 445148 239220 445176
rect 238812 445136 238818 445148
rect 239214 445136 239220 445148
rect 239272 445136 239278 445188
rect 240502 445136 240508 445188
rect 240560 445176 240566 445188
rect 241146 445176 241152 445188
rect 240560 445148 241152 445176
rect 240560 445136 240566 445148
rect 241146 445136 241152 445148
rect 241204 445136 241210 445188
rect 241790 445136 241796 445188
rect 241848 445176 241854 445188
rect 242434 445176 242440 445188
rect 241848 445148 242440 445176
rect 241848 445136 241854 445148
rect 242434 445136 242440 445148
rect 242492 445136 242498 445188
rect 243078 445136 243084 445188
rect 243136 445176 243142 445188
rect 243906 445176 243912 445188
rect 243136 445148 243912 445176
rect 243136 445136 243142 445148
rect 243906 445136 243912 445148
rect 243964 445136 243970 445188
rect 244366 445136 244372 445188
rect 244424 445176 244430 445188
rect 245562 445176 245568 445188
rect 244424 445148 245568 445176
rect 244424 445136 244430 445148
rect 245562 445136 245568 445148
rect 245620 445136 245626 445188
rect 247310 445136 247316 445188
rect 247368 445176 247374 445188
rect 248138 445176 248144 445188
rect 247368 445148 248144 445176
rect 247368 445136 247374 445148
rect 248138 445136 248144 445148
rect 248196 445136 248202 445188
rect 248414 445136 248420 445188
rect 248472 445176 248478 445188
rect 249058 445176 249064 445188
rect 248472 445148 249064 445176
rect 248472 445136 248478 445148
rect 249058 445136 249064 445148
rect 249116 445136 249122 445188
rect 251818 445136 251824 445188
rect 251876 445176 251882 445188
rect 293862 445176 293868 445188
rect 251876 445148 293868 445176
rect 251876 445136 251882 445148
rect 293862 445136 293868 445148
rect 293920 445136 293926 445188
rect 3970 445068 3976 445120
rect 4028 445108 4034 445120
rect 216582 445108 216588 445120
rect 4028 445080 216588 445108
rect 4028 445068 4034 445080
rect 216582 445068 216588 445080
rect 216640 445068 216646 445120
rect 216766 445068 216772 445120
rect 216824 445108 216830 445120
rect 217778 445108 217784 445120
rect 216824 445080 217784 445108
rect 216824 445068 216830 445080
rect 217778 445068 217784 445080
rect 217836 445068 217842 445120
rect 218606 445068 218612 445120
rect 218664 445108 218670 445120
rect 219250 445108 219256 445120
rect 218664 445080 219256 445108
rect 218664 445068 218670 445080
rect 219250 445068 219256 445080
rect 219308 445068 219314 445120
rect 220814 445068 220820 445120
rect 220872 445108 220878 445120
rect 221274 445108 221280 445120
rect 220872 445080 221280 445108
rect 220872 445068 220878 445080
rect 221274 445068 221280 445080
rect 221332 445068 221338 445120
rect 224218 445068 224224 445120
rect 224276 445108 224282 445120
rect 224678 445108 224684 445120
rect 224276 445080 224684 445108
rect 224276 445068 224282 445080
rect 224678 445068 224684 445080
rect 224736 445068 224742 445120
rect 238846 445068 238852 445120
rect 238904 445108 238910 445120
rect 239858 445108 239864 445120
rect 238904 445080 239864 445108
rect 238904 445068 238910 445080
rect 239858 445068 239864 445080
rect 239916 445068 239922 445120
rect 244090 445068 244096 445120
rect 244148 445108 244154 445120
rect 293678 445108 293684 445120
rect 244148 445080 293684 445108
rect 244148 445068 244154 445080
rect 293678 445068 293684 445080
rect 293736 445068 293742 445120
rect 3234 445000 3240 445052
rect 3292 445040 3298 445052
rect 219342 445040 219348 445052
rect 3292 445012 219348 445040
rect 3292 445000 3298 445012
rect 219342 445000 219348 445012
rect 219400 445000 219406 445052
rect 248598 445000 248604 445052
rect 248656 445040 248662 445052
rect 299474 445040 299480 445052
rect 248656 445012 299480 445040
rect 248656 445000 248662 445012
rect 299474 445000 299480 445012
rect 299532 445000 299538 445052
rect 212994 444932 213000 444984
rect 213052 444972 213058 444984
rect 265710 444972 265716 444984
rect 213052 444944 265716 444972
rect 213052 444932 213058 444944
rect 265710 444932 265716 444944
rect 265768 444932 265774 444984
rect 199470 444864 199476 444916
rect 199528 444904 199534 444916
rect 227346 444904 227352 444916
rect 199528 444876 227352 444904
rect 199528 444864 199534 444876
rect 227346 444864 227352 444876
rect 227404 444864 227410 444916
rect 240226 444864 240232 444916
rect 240284 444904 240290 444916
rect 293586 444904 293592 444916
rect 240284 444876 293592 444904
rect 240284 444864 240290 444876
rect 293586 444864 293592 444876
rect 293644 444864 293650 444916
rect 199378 444796 199384 444848
rect 199436 444836 199442 444848
rect 228450 444836 228456 444848
rect 199436 444808 228456 444836
rect 199436 444796 199442 444808
rect 228450 444796 228456 444808
rect 228508 444796 228514 444848
rect 235442 444796 235448 444848
rect 235500 444836 235506 444848
rect 293494 444836 293500 444848
rect 235500 444808 293500 444836
rect 235500 444796 235506 444808
rect 293494 444796 293500 444808
rect 293552 444796 293558 444848
rect 211890 444728 211896 444780
rect 211948 444768 211954 444780
rect 269850 444768 269856 444780
rect 211948 444740 269856 444768
rect 211948 444728 211954 444740
rect 269850 444728 269856 444740
rect 269908 444728 269914 444780
rect 211338 444660 211344 444712
rect 211396 444700 211402 444712
rect 211396 444672 220032 444700
rect 211396 444660 211402 444672
rect 217042 444592 217048 444644
rect 217100 444632 217106 444644
rect 217318 444632 217324 444644
rect 217100 444604 217324 444632
rect 217100 444592 217106 444604
rect 217318 444592 217324 444604
rect 217376 444592 217382 444644
rect 220004 444632 220032 444672
rect 220078 444660 220084 444712
rect 220136 444700 220142 444712
rect 271230 444700 271236 444712
rect 220136 444672 271236 444700
rect 220136 444660 220142 444672
rect 271230 444660 271236 444672
rect 271288 444660 271294 444712
rect 273990 444632 273996 444644
rect 219360 444604 219572 444632
rect 220004 444604 273996 444632
rect 196618 444524 196624 444576
rect 196676 444564 196682 444576
rect 219360 444564 219388 444604
rect 196676 444536 219388 444564
rect 219544 444564 219572 444604
rect 273990 444592 273996 444604
rect 274048 444592 274054 444644
rect 227898 444564 227904 444576
rect 219544 444536 227904 444564
rect 196676 444524 196682 444536
rect 227898 444524 227904 444536
rect 227956 444524 227962 444576
rect 230474 444524 230480 444576
rect 230532 444564 230538 444576
rect 298646 444564 298652 444576
rect 230532 444536 298652 444564
rect 230532 444524 230538 444536
rect 298646 444524 298652 444536
rect 298704 444524 298710 444576
rect 213914 444456 213920 444508
rect 213972 444496 213978 444508
rect 295886 444496 295892 444508
rect 213972 444468 295892 444496
rect 213972 444456 213978 444468
rect 295886 444456 295892 444468
rect 295944 444456 295950 444508
rect 200850 444388 200856 444440
rect 200908 444428 200914 444440
rect 229002 444428 229008 444440
rect 200908 444400 229008 444428
rect 200908 444388 200914 444400
rect 229002 444388 229008 444400
rect 229060 444428 229066 444440
rect 299842 444428 299848 444440
rect 229060 444400 299848 444428
rect 229060 444388 229066 444400
rect 299842 444388 299848 444400
rect 299900 444388 299906 444440
rect 255406 443980 255412 444032
rect 255464 444020 255470 444032
rect 295794 444020 295800 444032
rect 255464 443992 295800 444020
rect 255464 443980 255470 443992
rect 295794 443980 295800 443992
rect 295852 443980 295858 444032
rect 255590 443912 255596 443964
rect 255648 443952 255654 443964
rect 297450 443952 297456 443964
rect 255648 443924 297456 443952
rect 255648 443912 255654 443924
rect 297450 443912 297456 443924
rect 297508 443912 297514 443964
rect 226518 443844 226524 443896
rect 226576 443844 226582 443896
rect 254302 443844 254308 443896
rect 254360 443884 254366 443896
rect 297634 443884 297640 443896
rect 254360 443856 297640 443884
rect 254360 443844 254366 443856
rect 297634 443844 297640 443856
rect 297692 443844 297698 443896
rect 226536 443816 226564 443844
rect 215266 443788 226564 443816
rect 200942 443368 200948 443420
rect 201000 443408 201006 443420
rect 215266 443408 215294 443788
rect 252646 443776 252652 443828
rect 252704 443816 252710 443828
rect 296898 443816 296904 443828
rect 252704 443788 296904 443816
rect 252704 443776 252710 443788
rect 296898 443776 296904 443788
rect 296956 443776 296962 443828
rect 201000 443380 215294 443408
rect 217336 443720 220308 443748
rect 201000 443368 201006 443380
rect 200758 443300 200764 443352
rect 200816 443340 200822 443352
rect 217336 443340 217364 443720
rect 220280 443680 220308 443720
rect 220446 443708 220452 443760
rect 220504 443748 220510 443760
rect 229462 443748 229468 443760
rect 220504 443720 229468 443748
rect 220504 443708 220510 443720
rect 229462 443708 229468 443720
rect 229520 443708 229526 443760
rect 249886 443708 249892 443760
rect 249944 443748 249950 443760
rect 297358 443748 297364 443760
rect 249944 443720 297364 443748
rect 249944 443708 249950 443720
rect 297358 443708 297364 443720
rect 297416 443708 297422 443760
rect 229830 443680 229836 443692
rect 220280 443652 229836 443680
rect 229830 443640 229836 443652
rect 229888 443640 229894 443692
rect 245654 443640 245660 443692
rect 245712 443680 245718 443692
rect 297542 443680 297548 443692
rect 245712 443652 297548 443680
rect 245712 443640 245718 443652
rect 297542 443640 297548 443652
rect 297600 443640 297606 443692
rect 220446 443612 220452 443624
rect 200816 443312 217364 443340
rect 217428 443584 220452 443612
rect 200816 443300 200822 443312
rect 197998 443232 198004 443284
rect 198056 443272 198062 443284
rect 217428 443272 217456 443584
rect 220446 443572 220452 443584
rect 220504 443572 220510 443624
rect 228174 443544 228180 443556
rect 198056 443244 217456 443272
rect 220188 443516 228180 443544
rect 198056 443232 198062 443244
rect 192478 443164 192484 443216
rect 192536 443204 192542 443216
rect 220188 443204 220216 443516
rect 228174 443504 228180 443516
rect 228232 443504 228238 443556
rect 225782 443476 225788 443488
rect 192536 443176 220216 443204
rect 224926 443448 225788 443476
rect 192536 443164 192542 443176
rect 4062 443096 4068 443148
rect 4120 443136 4126 443148
rect 224926 443136 224954 443448
rect 225782 443436 225788 443448
rect 225840 443436 225846 443488
rect 231826 443448 243032 443476
rect 225230 443368 225236 443420
rect 225288 443368 225294 443420
rect 227990 443368 227996 443420
rect 228048 443368 228054 443420
rect 230382 443368 230388 443420
rect 230440 443368 230446 443420
rect 4120 443108 224954 443136
rect 4120 443096 4126 443108
rect 3326 443028 3332 443080
rect 3384 443068 3390 443080
rect 225248 443068 225276 443368
rect 3384 443040 225276 443068
rect 3384 443028 3390 443040
rect 3602 442960 3608 443012
rect 3660 443000 3666 443012
rect 228008 443000 228036 443368
rect 230400 443136 230428 443368
rect 231826 443136 231854 443448
rect 233694 443368 233700 443420
rect 233752 443408 233758 443420
rect 233752 443380 237420 443408
rect 233752 443368 233758 443380
rect 230400 443108 231854 443136
rect 3660 442972 228036 443000
rect 237392 443000 237420 443380
rect 242894 443368 242900 443420
rect 242952 443368 242958 443420
rect 242912 443068 242940 443368
rect 243004 443204 243032 443448
rect 249702 443368 249708 443420
rect 249760 443408 249766 443420
rect 249760 443380 258074 443408
rect 249760 443368 249766 443380
rect 258046 443204 258074 443380
rect 275462 443204 275468 443216
rect 243004 443176 253934 443204
rect 258046 443176 275468 443204
rect 253906 443136 253934 443176
rect 275462 443164 275468 443176
rect 275520 443164 275526 443216
rect 275370 443136 275376 443148
rect 253906 443108 275376 443136
rect 275370 443096 275376 443108
rect 275428 443096 275434 443148
rect 296806 443068 296812 443080
rect 242912 443040 296812 443068
rect 296806 443028 296812 443040
rect 296864 443028 296870 443080
rect 298002 443000 298008 443012
rect 237392 442972 298008 443000
rect 3660 442960 3666 442972
rect 298002 442960 298008 442972
rect 298060 442960 298066 443012
rect 265894 431876 265900 431928
rect 265952 431916 265958 431928
rect 298002 431916 298008 431928
rect 265952 431888 298008 431916
rect 265952 431876 265958 431888
rect 298002 431876 298008 431888
rect 298060 431876 298066 431928
rect 384298 431876 384304 431928
rect 384356 431916 384362 431928
rect 580166 431916 580172 431928
rect 384356 431888 580172 431916
rect 384356 431876 384362 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 266998 426368 267004 426420
rect 267056 426408 267062 426420
rect 298002 426408 298008 426420
rect 267056 426380 298008 426408
rect 267056 426368 267062 426380
rect 298002 426368 298008 426380
rect 298060 426368 298066 426420
rect 2774 410932 2780 410984
rect 2832 410972 2838 410984
rect 4982 410972 4988 410984
rect 2832 410944 4988 410972
rect 2832 410932 2838 410944
rect 4982 410932 4988 410944
rect 5040 410932 5046 410984
rect 265802 404268 265808 404320
rect 265860 404308 265866 404320
rect 298002 404308 298008 404320
rect 265860 404280 298008 404308
rect 265860 404268 265866 404280
rect 298002 404268 298008 404280
rect 298060 404268 298066 404320
rect 293862 401548 293868 401600
rect 293920 401588 293926 401600
rect 385034 401588 385040 401600
rect 293920 401560 385040 401588
rect 293920 401548 293926 401560
rect 385034 401548 385040 401560
rect 385092 401548 385098 401600
rect 297174 401344 297180 401396
rect 297232 401384 297238 401396
rect 297232 401356 313274 401384
rect 297232 401344 297238 401356
rect 313246 401316 313274 401356
rect 313246 401288 314654 401316
rect 314626 401248 314654 401288
rect 309244 401220 314240 401248
rect 314626 401220 327074 401248
rect 293402 401072 293408 401124
rect 293460 401112 293466 401124
rect 298002 401112 298008 401124
rect 293460 401084 298008 401112
rect 293460 401072 293466 401084
rect 298002 401072 298008 401084
rect 298060 401072 298066 401124
rect 298756 401084 303614 401112
rect 292942 401004 292948 401056
rect 293000 401044 293006 401056
rect 298756 401044 298784 401084
rect 293000 401016 298784 401044
rect 303586 401044 303614 401084
rect 303586 401016 308352 401044
rect 293000 401004 293006 401016
rect 293218 400936 293224 400988
rect 293276 400976 293282 400988
rect 297174 400976 297180 400988
rect 293276 400948 297180 400976
rect 293276 400936 293282 400948
rect 297174 400936 297180 400948
rect 297232 400936 297238 400988
rect 308324 400976 308352 401016
rect 309244 400976 309272 401220
rect 314212 401112 314240 401220
rect 314212 401084 317414 401112
rect 308324 400948 309272 400976
rect 293310 400868 293316 400920
rect 293368 400908 293374 400920
rect 317386 400908 317414 401084
rect 318766 400948 321784 400976
rect 318766 400908 318794 400948
rect 293368 400880 304994 400908
rect 317386 400880 318794 400908
rect 293368 400868 293374 400880
rect 299658 400732 299664 400784
rect 299716 400772 299722 400784
rect 299842 400772 299848 400784
rect 299716 400744 299848 400772
rect 299716 400732 299722 400744
rect 299842 400732 299848 400744
rect 299900 400732 299906 400784
rect 304966 400772 304994 400880
rect 314626 400812 318794 400840
rect 314626 400772 314654 400812
rect 304966 400744 314654 400772
rect 298002 400664 298008 400716
rect 298060 400704 298066 400716
rect 307570 400704 307576 400716
rect 298060 400676 307576 400704
rect 298060 400664 298066 400676
rect 307570 400664 307576 400676
rect 307628 400664 307634 400716
rect 318766 400636 318794 400812
rect 321756 400704 321784 400948
rect 324222 400704 324228 400716
rect 321756 400676 324228 400704
rect 324222 400664 324228 400676
rect 324280 400664 324286 400716
rect 327046 400704 327074 401220
rect 332502 400704 332508 400716
rect 327046 400676 332508 400704
rect 332502 400664 332508 400676
rect 332560 400664 332566 400716
rect 340966 400704 340972 400716
rect 336706 400676 340972 400704
rect 336706 400636 336734 400676
rect 340966 400664 340972 400676
rect 341024 400664 341030 400716
rect 318766 400608 336734 400636
rect 298554 400120 298560 400172
rect 298612 400160 298618 400172
rect 579982 400160 579988 400172
rect 298612 400132 579988 400160
rect 298612 400120 298618 400132
rect 579982 400120 579988 400132
rect 580040 400120 580046 400172
rect 252646 399780 252652 399832
rect 252704 399820 252710 399832
rect 253474 399820 253480 399832
rect 252704 399792 253480 399820
rect 252704 399780 252710 399792
rect 253474 399780 253480 399792
rect 253532 399780 253538 399832
rect 252646 399644 252652 399696
rect 252704 399684 252710 399696
rect 253198 399684 253204 399696
rect 252704 399656 253204 399684
rect 252704 399644 252710 399656
rect 253198 399644 253204 399656
rect 253256 399644 253262 399696
rect 253198 399508 253204 399560
rect 253256 399548 253262 399560
rect 253658 399548 253664 399560
rect 253256 399520 253664 399548
rect 253256 399508 253262 399520
rect 253658 399508 253664 399520
rect 253716 399508 253722 399560
rect 253106 399372 253112 399424
rect 253164 399412 253170 399424
rect 253658 399412 253664 399424
rect 253164 399384 253664 399412
rect 253164 399372 253170 399384
rect 253658 399372 253664 399384
rect 253716 399372 253722 399424
rect 205634 399100 205640 399152
rect 205692 399140 205698 399152
rect 210234 399140 210240 399152
rect 205692 399112 210240 399140
rect 205692 399100 205698 399112
rect 210234 399100 210240 399112
rect 210292 399100 210298 399152
rect 207658 399032 207664 399084
rect 207716 399072 207722 399084
rect 207716 399044 214696 399072
rect 207716 399032 207722 399044
rect 214668 399004 214696 399044
rect 216950 399032 216956 399084
rect 217008 399072 217014 399084
rect 217686 399072 217692 399084
rect 217008 399044 217692 399072
rect 217008 399032 217014 399044
rect 217686 399032 217692 399044
rect 217744 399032 217750 399084
rect 220814 399004 220820 399016
rect 214668 398976 220820 399004
rect 220814 398964 220820 398976
rect 220872 398964 220878 399016
rect 244366 398964 244372 399016
rect 244424 399004 244430 399016
rect 437474 399004 437480 399016
rect 244424 398976 437480 399004
rect 244424 398964 244430 398976
rect 437474 398964 437480 398976
rect 437532 398964 437538 399016
rect 209866 398896 209872 398948
rect 209924 398936 209930 398948
rect 226702 398936 226708 398948
rect 209924 398908 226708 398936
rect 209924 398896 209930 398908
rect 226702 398896 226708 398908
rect 226760 398896 226766 398948
rect 244826 398896 244832 398948
rect 244884 398936 244890 398948
rect 244884 398908 251174 398936
rect 244884 398896 244890 398908
rect 210234 398828 210240 398880
rect 210292 398868 210298 398880
rect 226334 398868 226340 398880
rect 210292 398840 226340 398868
rect 210292 398828 210298 398840
rect 226334 398828 226340 398840
rect 226392 398828 226398 398880
rect 245930 398828 245936 398880
rect 245988 398868 245994 398880
rect 245988 398840 250392 398868
rect 245988 398828 245994 398840
rect 206278 398760 206284 398812
rect 206336 398800 206342 398812
rect 219434 398800 219440 398812
rect 206336 398772 219440 398800
rect 206336 398760 206342 398772
rect 219434 398760 219440 398772
rect 219492 398760 219498 398812
rect 230842 398800 230848 398812
rect 229066 398772 230848 398800
rect 217686 398692 217692 398744
rect 217744 398732 217750 398744
rect 227714 398732 227720 398744
rect 217744 398704 227720 398732
rect 217744 398692 217750 398704
rect 227714 398692 227720 398704
rect 227772 398692 227778 398744
rect 207750 398624 207756 398676
rect 207808 398664 207814 398676
rect 223390 398664 223396 398676
rect 207808 398636 223396 398664
rect 207808 398624 207814 398636
rect 223390 398624 223396 398636
rect 223448 398624 223454 398676
rect 211890 398556 211896 398608
rect 211948 398596 211954 398608
rect 213546 398596 213552 398608
rect 211948 398568 213552 398596
rect 211948 398556 211954 398568
rect 213546 398556 213552 398568
rect 213604 398556 213610 398608
rect 208394 398488 208400 398540
rect 208452 398528 208458 398540
rect 226518 398528 226524 398540
rect 208452 398500 226524 398528
rect 208452 398488 208458 398500
rect 226518 398488 226524 398500
rect 226576 398488 226582 398540
rect 208026 398420 208032 398472
rect 208084 398460 208090 398472
rect 218882 398460 218888 398472
rect 208084 398432 218888 398460
rect 208084 398420 208090 398432
rect 218882 398420 218888 398432
rect 218940 398420 218946 398472
rect 207014 398352 207020 398404
rect 207072 398392 207078 398404
rect 226426 398392 226432 398404
rect 207072 398364 226432 398392
rect 207072 398352 207078 398364
rect 226426 398352 226432 398364
rect 226484 398352 226490 398404
rect 189074 398284 189080 398336
rect 189132 398324 189138 398336
rect 225046 398324 225052 398336
rect 189132 398296 225052 398324
rect 189132 398284 189138 398296
rect 225046 398284 225052 398296
rect 225104 398284 225110 398336
rect 171134 398216 171140 398268
rect 171192 398256 171198 398268
rect 223666 398256 223672 398268
rect 171192 398228 223672 398256
rect 171192 398216 171198 398228
rect 223666 398216 223672 398228
rect 223724 398216 223730 398268
rect 164234 398148 164240 398200
rect 164292 398188 164298 398200
rect 164292 398160 218744 398188
rect 164292 398148 164298 398160
rect 125594 398080 125600 398132
rect 125652 398120 125658 398132
rect 125652 398092 205634 398120
rect 125652 398080 125658 398092
rect 205606 397984 205634 398092
rect 211430 398080 211436 398132
rect 211488 398120 211494 398132
rect 212442 398120 212448 398132
rect 211488 398092 212448 398120
rect 211488 398080 211494 398092
rect 212442 398080 212448 398092
rect 212500 398080 212506 398132
rect 218606 398120 218612 398132
rect 215128 398092 218612 398120
rect 209314 398012 209320 398064
rect 209372 398052 209378 398064
rect 215128 398052 215156 398092
rect 218606 398080 218612 398092
rect 218664 398080 218670 398132
rect 209372 398024 215156 398052
rect 209372 398012 209378 398024
rect 212810 397984 212816 397996
rect 205606 397956 212816 397984
rect 212810 397944 212816 397956
rect 212868 397944 212874 397996
rect 218716 397984 218744 398160
rect 218882 398148 218888 398200
rect 218940 398188 218946 398200
rect 219342 398188 219348 398200
rect 218940 398160 219348 398188
rect 218940 398148 218946 398160
rect 219342 398148 219348 398160
rect 219400 398148 219406 398200
rect 219342 398012 219348 398064
rect 219400 398052 219406 398064
rect 229066 398052 229094 398772
rect 230842 398760 230848 398772
rect 230900 398760 230906 398812
rect 242618 398760 242624 398812
rect 242676 398800 242682 398812
rect 242676 398772 250208 398800
rect 242676 398760 242682 398772
rect 250180 398744 250208 398772
rect 250162 398692 250168 398744
rect 250220 398692 250226 398744
rect 250364 398596 250392 398840
rect 251146 398732 251174 398908
rect 253474 398896 253480 398948
rect 253532 398936 253538 398948
rect 543734 398936 543740 398948
rect 253532 398908 543740 398936
rect 253532 398896 253538 398908
rect 543734 398896 543740 398908
rect 543792 398896 543798 398948
rect 254302 398828 254308 398880
rect 254360 398868 254366 398880
rect 564434 398868 564440 398880
rect 254360 398840 564440 398868
rect 254360 398828 254366 398840
rect 564434 398828 564440 398840
rect 564492 398828 564498 398880
rect 252738 398760 252744 398812
rect 252796 398800 252802 398812
rect 253106 398800 253112 398812
rect 252796 398772 253112 398800
rect 252796 398760 252802 398772
rect 253106 398760 253112 398772
rect 253164 398760 253170 398812
rect 261478 398800 261484 398812
rect 253906 398772 261484 398800
rect 253906 398732 253934 398772
rect 261478 398760 261484 398772
rect 261536 398760 261542 398812
rect 293586 398760 293592 398812
rect 293644 398800 293650 398812
rect 303890 398800 303896 398812
rect 293644 398772 303896 398800
rect 293644 398760 293650 398772
rect 303890 398760 303896 398772
rect 303948 398760 303954 398812
rect 251146 398704 253934 398732
rect 299382 398692 299388 398744
rect 299440 398732 299446 398744
rect 370866 398732 370872 398744
rect 299440 398704 370872 398732
rect 299440 398692 299446 398704
rect 370866 398692 370872 398704
rect 370924 398692 370930 398744
rect 251146 398636 253934 398664
rect 251146 398596 251174 398636
rect 246684 398568 249472 398596
rect 250364 398568 251174 398596
rect 253906 398596 253934 398636
rect 293678 398624 293684 398676
rect 293736 398664 293742 398676
rect 362494 398664 362500 398676
rect 293736 398636 362500 398664
rect 293736 398624 293742 398636
rect 362494 398624 362500 398636
rect 362552 398624 362558 398676
rect 264238 398596 264244 398608
rect 253906 398568 264244 398596
rect 246206 398488 246212 398540
rect 246264 398528 246270 398540
rect 246684 398528 246712 398568
rect 246264 398500 246712 398528
rect 246264 398488 246270 398500
rect 246758 398420 246764 398472
rect 246816 398460 246822 398472
rect 246816 398432 248920 398460
rect 246816 398420 246822 398432
rect 248892 398392 248920 398432
rect 249444 398392 249472 398568
rect 264238 398556 264244 398568
rect 264296 398556 264302 398608
rect 293770 398556 293776 398608
rect 293828 398596 293834 398608
rect 357986 398596 357992 398608
rect 293828 398568 357992 398596
rect 293828 398556 293834 398568
rect 357986 398556 357992 398568
rect 358044 398556 358050 398608
rect 253474 398488 253480 398540
rect 253532 398528 253538 398540
rect 264330 398528 264336 398540
rect 253532 398500 264336 398528
rect 253532 398488 253538 398500
rect 264330 398488 264336 398500
rect 264388 398488 264394 398540
rect 295794 398488 295800 398540
rect 295852 398528 295858 398540
rect 354122 398528 354128 398540
rect 295852 398500 354128 398528
rect 295852 398488 295858 398500
rect 354122 398488 354128 398500
rect 354180 398488 354186 398540
rect 255406 398420 255412 398472
rect 255464 398460 255470 398472
rect 278038 398460 278044 398472
rect 255464 398432 278044 398460
rect 255464 398420 255470 398432
rect 278038 398420 278044 398432
rect 278096 398420 278102 398472
rect 293494 398420 293500 398472
rect 293552 398460 293558 398472
rect 349614 398460 349620 398472
rect 293552 398432 349620 398460
rect 293552 398420 293558 398432
rect 349614 398420 349620 398432
rect 349672 398420 349678 398472
rect 269758 398392 269764 398404
rect 248892 398364 249380 398392
rect 249444 398364 269764 398392
rect 247310 398284 247316 398336
rect 247368 398324 247374 398336
rect 249352 398324 249380 398364
rect 269758 398352 269764 398364
rect 269816 398352 269822 398404
rect 299658 398352 299664 398404
rect 299716 398392 299722 398404
rect 345750 398392 345756 398404
rect 299716 398364 345756 398392
rect 299716 398352 299722 398364
rect 345750 398352 345756 398364
rect 345808 398352 345814 398404
rect 271138 398324 271144 398336
rect 247368 398296 249288 398324
rect 249352 398296 271144 398324
rect 247368 398284 247374 398296
rect 249260 398256 249288 398296
rect 271138 398284 271144 398296
rect 271196 398284 271202 398336
rect 298646 398284 298652 398336
rect 298704 398324 298710 398336
rect 320634 398324 320640 398336
rect 298704 398296 320640 398324
rect 298704 398284 298710 398296
rect 320634 398284 320640 398296
rect 320692 398284 320698 398336
rect 274082 398256 274088 398268
rect 234586 398228 249196 398256
rect 249260 398228 274088 398256
rect 230290 398148 230296 398200
rect 230348 398188 230354 398200
rect 234586 398188 234614 398228
rect 230348 398160 234614 398188
rect 230348 398148 230354 398160
rect 241514 398148 241520 398200
rect 241572 398188 241578 398200
rect 248506 398188 248512 398200
rect 241572 398160 248512 398188
rect 241572 398148 241578 398160
rect 248506 398148 248512 398160
rect 248564 398148 248570 398200
rect 249168 398188 249196 398228
rect 274082 398216 274088 398228
rect 274140 398216 274146 398268
rect 275370 398216 275376 398268
rect 275428 398256 275434 398268
rect 312262 398256 312268 398268
rect 275428 398228 312268 398256
rect 275428 398216 275434 398228
rect 312262 398216 312268 398228
rect 312320 398216 312326 398268
rect 256694 398188 256700 398200
rect 249168 398160 256700 398188
rect 256694 398148 256700 398160
rect 256752 398148 256758 398200
rect 275462 398148 275468 398200
rect 275520 398188 275526 398200
rect 366358 398188 366364 398200
rect 275520 398160 366364 398188
rect 275520 398148 275526 398160
rect 366358 398148 366364 398160
rect 366416 398148 366422 398200
rect 238202 398080 238208 398132
rect 238260 398120 238266 398132
rect 246482 398120 246488 398132
rect 238260 398092 246488 398120
rect 238260 398080 238266 398092
rect 246482 398080 246488 398092
rect 246540 398080 246546 398132
rect 247678 398080 247684 398132
rect 247736 398120 247742 398132
rect 480254 398120 480260 398132
rect 247736 398092 480260 398120
rect 247736 398080 247742 398092
rect 480254 398080 480260 398092
rect 480312 398080 480318 398132
rect 219400 398024 229094 398052
rect 219400 398012 219406 398024
rect 233234 398012 233240 398064
rect 233292 398052 233298 398064
rect 241514 398052 241520 398064
rect 233292 398024 241520 398052
rect 233292 398012 233298 398024
rect 241514 398012 241520 398024
rect 241572 398012 241578 398064
rect 243722 398012 243728 398064
rect 243780 398052 243786 398064
rect 243780 398024 253934 398052
rect 243780 398012 243786 398024
rect 223114 397984 223120 397996
rect 218716 397956 223120 397984
rect 223114 397944 223120 397956
rect 223172 397944 223178 397996
rect 237374 397944 237380 397996
rect 237432 397984 237438 397996
rect 243906 397984 243912 397996
rect 237432 397956 243912 397984
rect 237432 397944 237438 397956
rect 243906 397944 243912 397956
rect 243964 397944 243970 397996
rect 245378 397944 245384 397996
rect 245436 397984 245442 397996
rect 253474 397984 253480 397996
rect 245436 397956 253480 397984
rect 245436 397944 245442 397956
rect 253474 397944 253480 397956
rect 253532 397944 253538 397996
rect 253906 397984 253934 398024
rect 255498 398012 255504 398064
rect 255556 398052 255562 398064
rect 258810 398052 258816 398064
rect 255556 398024 258816 398052
rect 255556 398012 255562 398024
rect 258810 398012 258816 398024
rect 258868 398012 258874 398064
rect 257522 397984 257528 397996
rect 253906 397956 257528 397984
rect 257522 397944 257528 397956
rect 257580 397944 257586 397996
rect 207842 397876 207848 397928
rect 207900 397916 207906 397928
rect 217778 397916 217784 397928
rect 207900 397888 217784 397916
rect 207900 397876 207906 397888
rect 217778 397876 217784 397888
rect 217836 397876 217842 397928
rect 239858 397876 239864 397928
rect 239916 397916 239922 397928
rect 242618 397916 242624 397928
rect 239916 397888 242624 397916
rect 239916 397876 239922 397888
rect 242618 397876 242624 397888
rect 242676 397876 242682 397928
rect 244274 397876 244280 397928
rect 244332 397916 244338 397928
rect 247310 397916 247316 397928
rect 244332 397888 247316 397916
rect 244332 397876 244338 397888
rect 247310 397876 247316 397888
rect 247368 397876 247374 397928
rect 207934 397808 207940 397860
rect 207992 397848 207998 397860
rect 207992 397820 215156 397848
rect 207992 397808 207998 397820
rect 215128 397780 215156 397820
rect 240502 397808 240508 397860
rect 240560 397848 240566 397860
rect 247954 397848 247960 397860
rect 240560 397820 247960 397848
rect 240560 397808 240566 397820
rect 247954 397808 247960 397820
rect 248012 397808 248018 397860
rect 248506 397808 248512 397860
rect 248564 397848 248570 397860
rect 248564 397820 248736 397848
rect 248564 397808 248570 397820
rect 218330 397780 218336 397792
rect 215128 397752 218336 397780
rect 218330 397740 218336 397752
rect 218388 397740 218394 397792
rect 222838 397780 222844 397792
rect 218440 397752 222844 397780
rect 209130 397672 209136 397724
rect 209188 397712 209194 397724
rect 212258 397712 212264 397724
rect 209188 397684 212264 397712
rect 209188 397672 209194 397684
rect 212258 397672 212264 397684
rect 212316 397672 212322 397724
rect 213914 397672 213920 397724
rect 213972 397712 213978 397724
rect 216398 397712 216404 397724
rect 213972 397684 216404 397712
rect 213972 397672 213978 397684
rect 216398 397672 216404 397684
rect 216456 397672 216462 397724
rect 217778 397672 217784 397724
rect 217836 397712 217842 397724
rect 218440 397712 218468 397752
rect 222838 397740 222844 397752
rect 222896 397740 222902 397792
rect 231946 397740 231952 397792
rect 232004 397780 232010 397792
rect 239858 397780 239864 397792
rect 232004 397752 239864 397780
rect 232004 397740 232010 397752
rect 239858 397740 239864 397752
rect 239916 397740 239922 397792
rect 240226 397740 240232 397792
rect 240284 397780 240290 397792
rect 247678 397780 247684 397792
rect 240284 397752 247684 397780
rect 240284 397740 240290 397752
rect 247678 397740 247684 397752
rect 247736 397740 247742 397792
rect 248708 397780 248736 397820
rect 250162 397808 250168 397860
rect 250220 397848 250226 397860
rect 257430 397848 257436 397860
rect 250220 397820 257436 397848
rect 250220 397808 250226 397820
rect 257430 397808 257436 397820
rect 257488 397808 257494 397860
rect 256326 397780 256332 397792
rect 248064 397752 248276 397780
rect 248708 397752 256332 397780
rect 217836 397684 218468 397712
rect 217836 397672 217842 397684
rect 219434 397672 219440 397724
rect 219492 397712 219498 397724
rect 227438 397712 227444 397724
rect 219492 397684 227444 397712
rect 219492 397672 219498 397684
rect 227438 397672 227444 397684
rect 227496 397672 227502 397724
rect 243170 397672 243176 397724
rect 243228 397712 243234 397724
rect 248064 397712 248092 397752
rect 243228 397684 248092 397712
rect 248248 397712 248276 397752
rect 256326 397740 256332 397752
rect 256384 397740 256390 397792
rect 255958 397712 255964 397724
rect 248248 397684 255964 397712
rect 243228 397672 243234 397684
rect 255958 397672 255964 397684
rect 256016 397672 256022 397724
rect 209222 397604 209228 397656
rect 209280 397644 209286 397656
rect 212166 397644 212172 397656
rect 209280 397616 212172 397644
rect 209280 397604 209286 397616
rect 212166 397604 212172 397616
rect 212224 397604 212230 397656
rect 213362 397604 213368 397656
rect 213420 397644 213426 397656
rect 217226 397644 217232 397656
rect 213420 397616 217232 397644
rect 213420 397604 213426 397616
rect 217226 397604 217232 397616
rect 217284 397604 217290 397656
rect 222194 397604 222200 397656
rect 222252 397644 222258 397656
rect 227622 397644 227628 397656
rect 222252 397616 227628 397644
rect 222252 397604 222258 397616
rect 227622 397604 227628 397616
rect 227680 397604 227686 397656
rect 234062 397604 234068 397656
rect 234120 397644 234126 397656
rect 234430 397644 234436 397656
rect 234120 397616 234436 397644
rect 234120 397604 234126 397616
rect 234430 397604 234436 397616
rect 234488 397604 234494 397656
rect 239306 397604 239312 397656
rect 239364 397644 239370 397656
rect 246942 397644 246948 397656
rect 239364 397616 246948 397644
rect 239364 397604 239370 397616
rect 246942 397604 246948 397616
rect 247000 397604 247006 397656
rect 247310 397604 247316 397656
rect 247368 397644 247374 397656
rect 258718 397644 258724 397656
rect 247368 397616 258724 397644
rect 247368 397604 247374 397616
rect 258718 397604 258724 397616
rect 258776 397604 258782 397656
rect 215018 397576 215024 397588
rect 212368 397548 215024 397576
rect 212166 397468 212172 397520
rect 212224 397508 212230 397520
rect 212368 397508 212396 397548
rect 215018 397536 215024 397548
rect 215076 397536 215082 397588
rect 216398 397536 216404 397588
rect 216456 397576 216462 397588
rect 222378 397576 222384 397588
rect 216456 397548 222384 397576
rect 216456 397536 216462 397548
rect 222378 397536 222384 397548
rect 222436 397536 222442 397588
rect 226334 397536 226340 397588
rect 226392 397576 226398 397588
rect 227898 397576 227904 397588
rect 226392 397548 227904 397576
rect 226392 397536 226398 397548
rect 227898 397536 227904 397548
rect 227956 397536 227962 397588
rect 242066 397536 242072 397588
rect 242124 397576 242130 397588
rect 256142 397576 256148 397588
rect 242124 397548 256148 397576
rect 242124 397536 242130 397548
rect 256142 397536 256148 397548
rect 256200 397536 256206 397588
rect 256234 397536 256240 397588
rect 256292 397576 256298 397588
rect 256292 397548 258074 397576
rect 256292 397536 256298 397548
rect 212224 397480 212396 397508
rect 212224 397468 212230 397480
rect 212810 397468 212816 397520
rect 212868 397508 212874 397520
rect 220078 397508 220084 397520
rect 212868 397480 220084 397508
rect 212868 397468 212874 397480
rect 220078 397468 220084 397480
rect 220136 397468 220142 397520
rect 227622 397468 227628 397520
rect 227680 397508 227686 397520
rect 228266 397508 228272 397520
rect 227680 397480 228272 397508
rect 227680 397468 227686 397480
rect 228266 397468 228272 397480
rect 228324 397468 228330 397520
rect 231486 397468 231492 397520
rect 231544 397508 231550 397520
rect 234062 397508 234068 397520
rect 231544 397480 234068 397508
rect 231544 397468 231550 397480
rect 234062 397468 234068 397480
rect 234120 397468 234126 397520
rect 236086 397468 236092 397520
rect 236144 397508 236150 397520
rect 238202 397508 238208 397520
rect 236144 397480 238208 397508
rect 236144 397468 236150 397480
rect 238202 397468 238208 397480
rect 238260 397468 238266 397520
rect 238754 397468 238760 397520
rect 238812 397508 238818 397520
rect 244826 397508 244832 397520
rect 238812 397480 244832 397508
rect 238812 397468 238818 397480
rect 244826 397468 244832 397480
rect 244884 397468 244890 397520
rect 258046 397508 258074 397548
rect 525794 397508 525800 397520
rect 258046 397480 525800 397508
rect 525794 397468 525800 397480
rect 525852 397468 525858 397520
rect 255958 397332 255964 397384
rect 256016 397372 256022 397384
rect 256142 397372 256148 397384
rect 256016 397344 256148 397372
rect 256016 397332 256022 397344
rect 256142 397332 256148 397344
rect 256200 397332 256206 397384
rect 201494 397264 201500 397316
rect 201552 397304 201558 397316
rect 226058 397304 226064 397316
rect 201552 397276 226064 397304
rect 201552 397264 201558 397276
rect 226058 397264 226064 397276
rect 226116 397264 226122 397316
rect 209038 397196 209044 397248
rect 209096 397236 209102 397248
rect 224678 397236 224684 397248
rect 209096 397208 224684 397236
rect 209096 397196 209102 397208
rect 224678 397196 224684 397208
rect 224736 397196 224742 397248
rect 194594 397128 194600 397180
rect 194652 397168 194658 397180
rect 225506 397168 225512 397180
rect 194652 397140 225512 397168
rect 194652 397128 194658 397140
rect 225506 397128 225512 397140
rect 225564 397128 225570 397180
rect 237006 397128 237012 397180
rect 237064 397168 237070 397180
rect 237064 397140 244274 397168
rect 237064 397128 237070 397140
rect 155954 397060 155960 397112
rect 156012 397100 156018 397112
rect 222470 397100 222476 397112
rect 156012 397072 222476 397100
rect 156012 397060 156018 397072
rect 222470 397060 222476 397072
rect 222528 397060 222534 397112
rect 225598 397060 225604 397112
rect 225656 397100 225662 397112
rect 226058 397100 226064 397112
rect 225656 397072 226064 397100
rect 225656 397060 225662 397072
rect 226058 397060 226064 397072
rect 226116 397060 226122 397112
rect 230474 397060 230480 397112
rect 230532 397100 230538 397112
rect 242066 397100 242072 397112
rect 230532 397072 242072 397100
rect 230532 397060 230538 397072
rect 242066 397060 242072 397072
rect 242124 397060 242130 397112
rect 244246 397100 244274 397140
rect 251542 397128 251548 397180
rect 251600 397168 251606 397180
rect 255958 397168 255964 397180
rect 251600 397140 255964 397168
rect 251600 397128 251606 397140
rect 255958 397128 255964 397140
rect 256016 397128 256022 397180
rect 244246 397072 253934 397100
rect 144914 396992 144920 397044
rect 144972 397032 144978 397044
rect 221642 397032 221648 397044
rect 144972 397004 221648 397032
rect 144972 396992 144978 397004
rect 221642 396992 221648 397004
rect 221700 396992 221706 397044
rect 229186 396992 229192 397044
rect 229244 397032 229250 397044
rect 230198 397032 230204 397044
rect 229244 397004 230204 397032
rect 229244 396992 229250 397004
rect 230198 396992 230204 397004
rect 230256 396992 230262 397044
rect 232682 396992 232688 397044
rect 232740 397032 232746 397044
rect 232866 397032 232872 397044
rect 232740 397004 232872 397032
rect 232740 396992 232746 397004
rect 232866 396992 232872 397004
rect 232924 396992 232930 397044
rect 241698 396992 241704 397044
rect 241756 397032 241762 397044
rect 241756 397004 249104 397032
rect 241756 396992 241762 397004
rect 131114 396924 131120 396976
rect 131172 396964 131178 396976
rect 131172 396936 214052 396964
rect 131172 396924 131178 396936
rect 77294 396856 77300 396908
rect 77352 396896 77358 396908
rect 213914 396896 213920 396908
rect 77352 396868 213920 396896
rect 77352 396856 77358 396868
rect 213914 396856 213920 396868
rect 213972 396856 213978 396908
rect 46934 396788 46940 396840
rect 46992 396828 46998 396840
rect 211154 396828 211160 396840
rect 46992 396800 211160 396828
rect 46992 396788 46998 396800
rect 211154 396788 211160 396800
rect 211212 396788 211218 396840
rect 214024 396828 214052 396936
rect 227806 396924 227812 396976
rect 227864 396964 227870 396976
rect 228634 396964 228640 396976
rect 227864 396936 228640 396964
rect 227864 396924 227870 396936
rect 228634 396924 228640 396936
rect 228692 396924 228698 396976
rect 229278 396924 229284 396976
rect 229336 396964 229342 396976
rect 230106 396964 230112 396976
rect 229336 396936 230112 396964
rect 229336 396924 229342 396936
rect 230106 396924 230112 396936
rect 230164 396924 230170 396976
rect 231854 396924 231860 396976
rect 231912 396964 231918 396976
rect 232958 396964 232964 396976
rect 231912 396936 232964 396964
rect 231912 396924 231918 396936
rect 232958 396924 232964 396936
rect 233016 396924 233022 396976
rect 225322 396856 225328 396908
rect 225380 396896 225386 396908
rect 225874 396896 225880 396908
rect 225380 396868 225880 396896
rect 225380 396856 225386 396868
rect 225874 396856 225880 396868
rect 225932 396856 225938 396908
rect 229370 396856 229376 396908
rect 229428 396896 229434 396908
rect 230014 396896 230020 396908
rect 229428 396868 230020 396896
rect 229428 396856 229434 396868
rect 230014 396856 230020 396868
rect 230072 396856 230078 396908
rect 231026 396856 231032 396908
rect 231084 396896 231090 396908
rect 231486 396896 231492 396908
rect 231084 396868 231492 396896
rect 231084 396856 231090 396868
rect 231486 396856 231492 396868
rect 231544 396856 231550 396908
rect 249076 396896 249104 397004
rect 253906 396964 253934 397072
rect 254210 396992 254216 397044
rect 254268 397032 254274 397044
rect 255038 397032 255044 397044
rect 254268 397004 255044 397032
rect 254268 396992 254274 397004
rect 255038 396992 255044 397004
rect 255096 396992 255102 397044
rect 342254 396964 342260 396976
rect 253906 396936 342260 396964
rect 342254 396924 342260 396936
rect 342312 396924 342318 396976
rect 402974 396896 402980 396908
rect 249076 396868 402980 396896
rect 402974 396856 402980 396868
rect 403032 396856 403038 396908
rect 220538 396828 220544 396840
rect 214024 396800 220544 396828
rect 220538 396788 220544 396800
rect 220596 396788 220602 396840
rect 228082 396788 228088 396840
rect 228140 396828 228146 396840
rect 228634 396828 228640 396840
rect 228140 396800 228640 396828
rect 228140 396788 228146 396800
rect 228634 396788 228640 396800
rect 228692 396788 228698 396840
rect 230566 396788 230572 396840
rect 230624 396828 230630 396840
rect 231762 396828 231768 396840
rect 230624 396800 231768 396828
rect 230624 396788 230630 396800
rect 231762 396788 231768 396800
rect 231820 396788 231826 396840
rect 231854 396788 231860 396840
rect 231912 396828 231918 396840
rect 232314 396828 232320 396840
rect 231912 396800 232320 396828
rect 231912 396788 231918 396800
rect 232314 396788 232320 396800
rect 232372 396788 232378 396840
rect 233602 396788 233608 396840
rect 233660 396828 233666 396840
rect 234246 396828 234252 396840
rect 233660 396800 234252 396828
rect 233660 396788 233666 396800
rect 234246 396788 234252 396800
rect 234304 396788 234310 396840
rect 242250 396788 242256 396840
rect 242308 396828 242314 396840
rect 409874 396828 409880 396840
rect 242308 396800 409880 396828
rect 242308 396788 242314 396800
rect 409874 396788 409880 396800
rect 409932 396788 409938 396840
rect 40034 396720 40040 396772
rect 40092 396760 40098 396772
rect 40092 396732 205634 396760
rect 40092 396720 40098 396732
rect 205606 396692 205634 396732
rect 226610 396720 226616 396772
rect 226668 396760 226674 396772
rect 227254 396760 227260 396772
rect 226668 396732 227260 396760
rect 226668 396720 226674 396732
rect 227254 396720 227260 396732
rect 227312 396720 227318 396772
rect 229738 396760 229744 396772
rect 229296 396732 229744 396760
rect 229296 396704 229324 396732
rect 229738 396720 229744 396732
rect 229796 396720 229802 396772
rect 230750 396720 230756 396772
rect 230808 396760 230814 396772
rect 231026 396760 231032 396772
rect 230808 396732 231032 396760
rect 230808 396720 230814 396732
rect 231026 396720 231032 396732
rect 231084 396720 231090 396772
rect 232222 396720 232228 396772
rect 232280 396760 232286 396772
rect 232590 396760 232596 396772
rect 232280 396732 232596 396760
rect 232280 396720 232286 396732
rect 232590 396720 232596 396732
rect 232648 396720 232654 396772
rect 233510 396720 233516 396772
rect 233568 396760 233574 396772
rect 233878 396760 233884 396772
rect 233568 396732 233884 396760
rect 233568 396720 233574 396732
rect 233878 396720 233884 396732
rect 233936 396720 233942 396772
rect 247218 396720 247224 396772
rect 247276 396760 247282 396772
rect 473354 396760 473360 396772
rect 247276 396732 473360 396760
rect 247276 396720 247282 396732
rect 473354 396720 473360 396732
rect 473412 396720 473418 396772
rect 213454 396692 213460 396704
rect 205606 396664 213460 396692
rect 213454 396652 213460 396664
rect 213512 396652 213518 396704
rect 225138 396652 225144 396704
rect 225196 396692 225202 396704
rect 226242 396692 226248 396704
rect 225196 396664 226248 396692
rect 225196 396652 225202 396664
rect 226242 396652 226248 396664
rect 226300 396652 226306 396704
rect 226702 396652 226708 396704
rect 226760 396692 226766 396704
rect 227162 396692 227168 396704
rect 226760 396664 227168 396692
rect 226760 396652 226766 396664
rect 227162 396652 227168 396664
rect 227220 396652 227226 396704
rect 229278 396652 229284 396704
rect 229336 396652 229342 396704
rect 230566 396652 230572 396704
rect 230624 396692 230630 396704
rect 231394 396692 231400 396704
rect 230624 396664 231400 396692
rect 230624 396652 230630 396664
rect 231394 396652 231400 396664
rect 231452 396652 231458 396704
rect 254026 396652 254032 396704
rect 254084 396692 254090 396704
rect 254854 396692 254860 396704
rect 254084 396664 254860 396692
rect 254084 396652 254090 396664
rect 254854 396652 254860 396664
rect 254912 396652 254918 396704
rect 225782 396584 225788 396636
rect 225840 396624 225846 396636
rect 225966 396624 225972 396636
rect 225840 396596 225972 396624
rect 225840 396584 225846 396596
rect 225966 396584 225972 396596
rect 226024 396584 226030 396636
rect 226518 396584 226524 396636
rect 226576 396624 226582 396636
rect 226978 396624 226984 396636
rect 226576 396596 226984 396624
rect 226576 396584 226582 396596
rect 226978 396584 226984 396596
rect 227036 396584 227042 396636
rect 225598 396516 225604 396568
rect 225656 396556 225662 396568
rect 227070 396556 227076 396568
rect 225656 396528 227076 396556
rect 225656 396516 225662 396528
rect 227070 396516 227076 396528
rect 227128 396516 227134 396568
rect 229094 396516 229100 396568
rect 229152 396556 229158 396568
rect 229462 396556 229468 396568
rect 229152 396528 229468 396556
rect 229152 396516 229158 396528
rect 229462 396516 229468 396528
rect 229520 396516 229526 396568
rect 229646 396516 229652 396568
rect 229704 396556 229710 396568
rect 229830 396556 229836 396568
rect 229704 396528 229836 396556
rect 229704 396516 229710 396528
rect 229830 396516 229836 396528
rect 229888 396516 229894 396568
rect 230750 396516 230756 396568
rect 230808 396556 230814 396568
rect 231118 396556 231124 396568
rect 230808 396528 231124 396556
rect 230808 396516 230814 396528
rect 231118 396516 231124 396528
rect 231176 396516 231182 396568
rect 232038 396516 232044 396568
rect 232096 396556 232102 396568
rect 232682 396556 232688 396568
rect 232096 396528 232688 396556
rect 232096 396516 232102 396528
rect 232682 396516 232688 396528
rect 232740 396516 232746 396568
rect 233510 396516 233516 396568
rect 233568 396556 233574 396568
rect 233970 396556 233976 396568
rect 233568 396528 233976 396556
rect 233568 396516 233574 396528
rect 233970 396516 233976 396528
rect 234028 396516 234034 396568
rect 254118 396516 254124 396568
rect 254176 396556 254182 396568
rect 254394 396556 254400 396568
rect 254176 396528 254400 396556
rect 254176 396516 254182 396528
rect 254394 396516 254400 396528
rect 254452 396516 254458 396568
rect 227990 396448 227996 396500
rect 228048 396448 228054 396500
rect 230658 396448 230664 396500
rect 230716 396488 230722 396500
rect 231210 396488 231216 396500
rect 230716 396460 231216 396488
rect 230716 396448 230722 396460
rect 231210 396448 231216 396460
rect 231268 396448 231274 396500
rect 232130 396448 232136 396500
rect 232188 396488 232194 396500
rect 232866 396488 232872 396500
rect 232188 396460 232872 396488
rect 232188 396448 232194 396460
rect 232866 396448 232872 396460
rect 232924 396448 232930 396500
rect 233418 396448 233424 396500
rect 233476 396488 233482 396500
rect 234154 396488 234160 396500
rect 233476 396460 234160 396488
rect 233476 396448 233482 396460
rect 234154 396448 234160 396460
rect 234212 396448 234218 396500
rect 226886 396244 226892 396296
rect 226944 396284 226950 396296
rect 227530 396284 227536 396296
rect 226944 396256 227536 396284
rect 226944 396244 226950 396256
rect 227530 396244 227536 396256
rect 227588 396244 227594 396296
rect 228008 396284 228036 396448
rect 234522 396380 234528 396432
rect 234580 396420 234586 396432
rect 235442 396420 235448 396432
rect 234580 396392 235448 396420
rect 234580 396380 234586 396392
rect 235442 396380 235448 396392
rect 235500 396380 235506 396432
rect 254302 396380 254308 396432
rect 254360 396420 254366 396432
rect 254670 396420 254676 396432
rect 254360 396392 254676 396420
rect 254360 396380 254366 396392
rect 254670 396380 254676 396392
rect 254728 396380 254734 396432
rect 254118 396312 254124 396364
rect 254176 396352 254182 396364
rect 254578 396352 254584 396364
rect 254176 396324 254584 396352
rect 254176 396312 254182 396324
rect 254578 396312 254584 396324
rect 254636 396312 254642 396364
rect 228174 396284 228180 396296
rect 228008 396256 228180 396284
rect 228174 396244 228180 396256
rect 228232 396244 228238 396296
rect 233878 396244 233884 396296
rect 233936 396284 233942 396296
rect 234062 396284 234068 396296
rect 233936 396256 234068 396284
rect 233936 396244 233942 396256
rect 234062 396244 234068 396256
rect 234120 396244 234126 396296
rect 253934 396108 253940 396160
rect 253992 396148 253998 396160
rect 254946 396148 254952 396160
rect 253992 396120 254952 396148
rect 253992 396108 253998 396120
rect 254946 396108 254952 396120
rect 255004 396108 255010 396160
rect 241606 395836 241612 395888
rect 241664 395876 241670 395888
rect 242434 395876 242440 395888
rect 241664 395848 242440 395876
rect 241664 395836 241670 395848
rect 242434 395836 242440 395848
rect 242492 395836 242498 395888
rect 248506 395836 248512 395888
rect 248564 395876 248570 395888
rect 249150 395876 249156 395888
rect 248564 395848 249156 395876
rect 248564 395836 248570 395848
rect 249150 395836 249156 395848
rect 249208 395836 249214 395888
rect 249242 395836 249248 395888
rect 249300 395876 249306 395888
rect 249518 395876 249524 395888
rect 249300 395848 249524 395876
rect 249300 395836 249306 395848
rect 249518 395836 249524 395848
rect 249576 395836 249582 395888
rect 231486 395768 231492 395820
rect 231544 395808 231550 395820
rect 266354 395808 266360 395820
rect 231544 395780 266360 395808
rect 231544 395768 231550 395780
rect 266354 395768 266360 395780
rect 266412 395768 266418 395820
rect 231302 395700 231308 395752
rect 231360 395740 231366 395752
rect 269114 395740 269120 395752
rect 231360 395712 269120 395740
rect 231360 395700 231366 395712
rect 269114 395700 269120 395712
rect 269172 395700 269178 395752
rect 232958 395632 232964 395684
rect 233016 395672 233022 395684
rect 276014 395672 276020 395684
rect 233016 395644 276020 395672
rect 233016 395632 233022 395644
rect 276014 395632 276020 395644
rect 276072 395632 276078 395684
rect 149698 395564 149704 395616
rect 149756 395604 149762 395616
rect 216950 395604 216956 395616
rect 149756 395576 216956 395604
rect 149756 395564 149762 395576
rect 216950 395564 216956 395576
rect 217008 395564 217014 395616
rect 241514 395564 241520 395616
rect 241572 395604 241578 395616
rect 293954 395604 293960 395616
rect 241572 395576 293960 395604
rect 241572 395564 241578 395576
rect 293954 395564 293960 395576
rect 294012 395564 294018 395616
rect 115934 395496 115940 395548
rect 115992 395536 115998 395548
rect 218882 395536 218888 395548
rect 115992 395508 218888 395536
rect 115992 395496 115998 395508
rect 218882 395496 218888 395508
rect 218940 395496 218946 395548
rect 223114 395496 223120 395548
rect 223172 395536 223178 395548
rect 227346 395536 227352 395548
rect 223172 395508 227352 395536
rect 223172 395496 223178 395508
rect 227346 395496 227352 395508
rect 227404 395496 227410 395548
rect 252002 395496 252008 395548
rect 252060 395536 252066 395548
rect 535454 395536 535460 395548
rect 252060 395508 535460 395536
rect 252060 395496 252066 395508
rect 535454 395496 535460 395508
rect 535512 395496 535518 395548
rect 52454 395428 52460 395480
rect 52512 395468 52518 395480
rect 214466 395468 214472 395480
rect 52512 395440 214472 395468
rect 52512 395428 52518 395440
rect 214466 395428 214472 395440
rect 214524 395428 214530 395480
rect 252646 395428 252652 395480
rect 252704 395468 252710 395480
rect 542354 395468 542360 395480
rect 252704 395440 542360 395468
rect 252704 395428 252710 395440
rect 542354 395428 542360 395440
rect 542412 395428 542418 395480
rect 30374 395360 30380 395412
rect 30432 395400 30438 395412
rect 212718 395400 212724 395412
rect 30432 395372 212724 395400
rect 30432 395360 30438 395372
rect 212718 395360 212724 395372
rect 212776 395360 212782 395412
rect 228358 395360 228364 395412
rect 228416 395400 228422 395412
rect 228542 395400 228548 395412
rect 228416 395372 228548 395400
rect 228416 395360 228422 395372
rect 228542 395360 228548 395372
rect 228600 395360 228606 395412
rect 253658 395360 253664 395412
rect 253716 395400 253722 395412
rect 549254 395400 549260 395412
rect 253716 395372 549260 395400
rect 253716 395360 253722 395372
rect 549254 395360 549260 395372
rect 549312 395360 549318 395412
rect 27614 395292 27620 395344
rect 27672 395332 27678 395344
rect 211430 395332 211436 395344
rect 27672 395304 211436 395332
rect 27672 395292 27678 395304
rect 211430 395292 211436 395304
rect 211488 395292 211494 395344
rect 255038 395292 255044 395344
rect 255096 395332 255102 395344
rect 564526 395332 564532 395344
rect 255096 395304 564532 395332
rect 255096 395292 255102 395304
rect 564526 395292 564532 395304
rect 564584 395292 564590 395344
rect 238846 395156 238852 395208
rect 238904 395196 238910 395208
rect 239766 395196 239772 395208
rect 238904 395168 239772 395196
rect 238904 395156 238910 395168
rect 239766 395156 239772 395168
rect 239824 395156 239830 395208
rect 244642 395088 244648 395140
rect 244700 395128 244706 395140
rect 245378 395128 245384 395140
rect 244700 395100 245384 395128
rect 244700 395088 244706 395100
rect 245378 395088 245384 395100
rect 245436 395088 245442 395140
rect 228266 394680 228272 394732
rect 228324 394720 228330 394732
rect 231118 394720 231124 394732
rect 228324 394692 231124 394720
rect 228324 394680 228330 394692
rect 231118 394680 231124 394692
rect 231176 394680 231182 394732
rect 232406 394680 232412 394732
rect 232464 394720 232470 394732
rect 232774 394720 232780 394732
rect 232464 394692 232780 394720
rect 232464 394680 232470 394692
rect 232774 394680 232780 394692
rect 232832 394680 232838 394732
rect 237926 394680 237932 394732
rect 237984 394720 237990 394732
rect 238386 394720 238392 394732
rect 237984 394692 238392 394720
rect 237984 394680 237990 394692
rect 238386 394680 238392 394692
rect 238444 394680 238450 394732
rect 235994 394612 236000 394664
rect 236052 394652 236058 394664
rect 243998 394652 244004 394664
rect 236052 394624 244004 394652
rect 236052 394612 236058 394624
rect 243998 394612 244004 394624
rect 244056 394612 244062 394664
rect 225230 394544 225236 394596
rect 225288 394584 225294 394596
rect 227714 394584 227720 394596
rect 225288 394556 227720 394584
rect 225288 394544 225294 394556
rect 227714 394544 227720 394556
rect 227772 394544 227778 394596
rect 228266 394544 228272 394596
rect 228324 394584 228330 394596
rect 228818 394584 228824 394596
rect 228324 394556 228824 394584
rect 228324 394544 228330 394556
rect 228818 394544 228824 394556
rect 228876 394544 228882 394596
rect 237374 394544 237380 394596
rect 237432 394584 237438 394596
rect 238018 394584 238024 394596
rect 237432 394556 238024 394584
rect 237432 394544 237438 394556
rect 238018 394544 238024 394556
rect 238076 394544 238082 394596
rect 251266 394544 251272 394596
rect 251324 394584 251330 394596
rect 251634 394584 251640 394596
rect 251324 394556 251640 394584
rect 251324 394544 251330 394556
rect 251634 394544 251640 394556
rect 251692 394544 251698 394596
rect 215294 394476 215300 394528
rect 215352 394516 215358 394528
rect 224218 394516 224224 394528
rect 215352 394488 224224 394516
rect 215352 394476 215358 394488
rect 224218 394476 224224 394488
rect 224276 394476 224282 394528
rect 234430 394476 234436 394528
rect 234488 394516 234494 394528
rect 304994 394516 305000 394528
rect 234488 394488 305000 394516
rect 234488 394476 234494 394488
rect 304994 394476 305000 394488
rect 305052 394476 305058 394528
rect 226150 394448 226156 394460
rect 215266 394420 226156 394448
rect 211982 394340 211988 394392
rect 212040 394380 212046 394392
rect 212534 394380 212540 394392
rect 212040 394352 212540 394380
rect 212040 394340 212046 394352
rect 212534 394340 212540 394352
rect 212592 394340 212598 394392
rect 214282 394340 214288 394392
rect 214340 394380 214346 394392
rect 214650 394380 214656 394392
rect 214340 394352 214656 394380
rect 214340 394340 214346 394352
rect 214650 394340 214656 394352
rect 214708 394340 214714 394392
rect 202874 394272 202880 394324
rect 202932 394312 202938 394324
rect 215266 394312 215294 394420
rect 226150 394408 226156 394420
rect 226208 394408 226214 394460
rect 235534 394408 235540 394460
rect 235592 394448 235598 394460
rect 235592 394420 237972 394448
rect 235592 394408 235598 394420
rect 234706 394340 234712 394392
rect 234764 394380 234770 394392
rect 235258 394380 235264 394392
rect 234764 394352 235264 394380
rect 234764 394340 234770 394352
rect 235258 394340 235264 394352
rect 235316 394340 235322 394392
rect 236270 394340 236276 394392
rect 236328 394380 236334 394392
rect 237944 394380 237972 394420
rect 238754 394408 238760 394460
rect 238812 394448 238818 394460
rect 239122 394448 239128 394460
rect 238812 394420 239128 394448
rect 238812 394408 238818 394420
rect 239122 394408 239128 394420
rect 239180 394408 239186 394460
rect 322934 394448 322940 394460
rect 239324 394420 322940 394448
rect 239324 394380 239352 394420
rect 322934 394408 322940 394420
rect 322992 394408 322998 394460
rect 236328 394352 237880 394380
rect 237944 394352 239352 394380
rect 239508 394352 241468 394380
rect 236328 394340 236334 394352
rect 202932 394284 215294 394312
rect 202932 394272 202938 394284
rect 221274 394272 221280 394324
rect 221332 394312 221338 394324
rect 221642 394312 221648 394324
rect 221332 394284 221648 394312
rect 221332 394272 221338 394284
rect 221642 394272 221648 394284
rect 221700 394272 221706 394324
rect 225046 394312 225052 394324
rect 224926 394284 225052 394312
rect 193214 394204 193220 394256
rect 193272 394244 193278 394256
rect 224926 394244 224954 394284
rect 225046 394272 225052 394284
rect 225104 394272 225110 394324
rect 193272 394216 224954 394244
rect 193272 394204 193278 394216
rect 229554 394204 229560 394256
rect 229612 394244 229618 394256
rect 229922 394244 229928 394256
rect 229612 394216 229928 394244
rect 229612 394204 229618 394216
rect 229922 394204 229928 394216
rect 229980 394204 229986 394256
rect 230198 394204 230204 394256
rect 230256 394244 230262 394256
rect 230256 394216 234614 394244
rect 230256 394204 230262 394216
rect 178034 394136 178040 394188
rect 178092 394176 178098 394188
rect 215294 394176 215300 394188
rect 178092 394148 215300 394176
rect 178092 394136 178098 394148
rect 215294 394136 215300 394148
rect 215352 394136 215358 394188
rect 220446 394176 220452 394188
rect 215404 394148 220452 394176
rect 129734 394068 129740 394120
rect 129792 394108 129798 394120
rect 215404 394108 215432 394148
rect 220446 394136 220452 394148
rect 220504 394136 220510 394188
rect 220998 394136 221004 394188
rect 221056 394176 221062 394188
rect 221458 394176 221464 394188
rect 221056 394148 221464 394176
rect 221056 394136 221062 394148
rect 221458 394136 221464 394148
rect 221516 394136 221522 394188
rect 234586 394176 234614 394216
rect 234890 394204 234896 394256
rect 234948 394244 234954 394256
rect 235258 394244 235264 394256
rect 234948 394216 235264 394244
rect 234948 394204 234954 394216
rect 235258 394204 235264 394216
rect 235316 394204 235322 394256
rect 237742 394244 237748 394256
rect 237576 394216 237748 394244
rect 236730 394176 236736 394188
rect 234586 394148 236736 394176
rect 236730 394136 236736 394148
rect 236788 394136 236794 394188
rect 215662 394108 215668 394120
rect 129792 394080 215432 394108
rect 215496 394080 215668 394108
rect 129792 394068 129798 394080
rect 69014 394000 69020 394052
rect 69072 394040 69078 394052
rect 215496 394040 215524 394080
rect 215662 394068 215668 394080
rect 215720 394068 215726 394120
rect 217042 394068 217048 394120
rect 217100 394108 217106 394120
rect 217410 394108 217416 394120
rect 217100 394080 217416 394108
rect 217100 394068 217106 394080
rect 217410 394068 217416 394080
rect 217468 394068 217474 394120
rect 219526 394068 219532 394120
rect 219584 394108 219590 394120
rect 220354 394108 220360 394120
rect 219584 394080 220360 394108
rect 219584 394068 219590 394080
rect 220354 394068 220360 394080
rect 220412 394068 220418 394120
rect 221182 394068 221188 394120
rect 221240 394108 221246 394120
rect 221550 394108 221556 394120
rect 221240 394080 221556 394108
rect 221240 394068 221246 394080
rect 221550 394068 221556 394080
rect 221608 394068 221614 394120
rect 234614 394068 234620 394120
rect 234672 394108 234678 394120
rect 234982 394108 234988 394120
rect 234672 394080 234988 394108
rect 234672 394068 234678 394080
rect 234982 394068 234988 394080
rect 235040 394068 235046 394120
rect 69072 394012 215524 394040
rect 69072 394000 69078 394012
rect 215570 394000 215576 394052
rect 215628 394040 215634 394052
rect 216306 394040 216312 394052
rect 215628 394012 216312 394040
rect 215628 394000 215634 394012
rect 216306 394000 216312 394012
rect 216364 394000 216370 394052
rect 216950 394000 216956 394052
rect 217008 394040 217014 394052
rect 217962 394040 217968 394052
rect 217008 394012 217968 394040
rect 217008 394000 217014 394012
rect 217962 394000 217968 394012
rect 218020 394000 218026 394052
rect 219618 394000 219624 394052
rect 219676 394040 219682 394052
rect 220170 394040 220176 394052
rect 219676 394012 220176 394040
rect 219676 394000 219682 394012
rect 220170 394000 220176 394012
rect 220228 394000 220234 394052
rect 220906 394000 220912 394052
rect 220964 394040 220970 394052
rect 221734 394040 221740 394052
rect 220964 394012 221740 394040
rect 220964 394000 220970 394012
rect 221734 394000 221740 394012
rect 221792 394000 221798 394052
rect 222378 394000 222384 394052
rect 222436 394040 222442 394052
rect 223206 394040 223212 394052
rect 222436 394012 223212 394040
rect 222436 394000 222442 394012
rect 223206 394000 223212 394012
rect 223264 394000 223270 394052
rect 223666 394000 223672 394052
rect 223724 394040 223730 394052
rect 224494 394040 224500 394052
rect 223724 394012 224500 394040
rect 223724 394000 223730 394012
rect 224494 394000 224500 394012
rect 224552 394000 224558 394052
rect 236086 394000 236092 394052
rect 236144 394040 236150 394052
rect 236362 394040 236368 394052
rect 236144 394012 236368 394040
rect 236144 394000 236150 394012
rect 236362 394000 236368 394012
rect 236420 394000 236426 394052
rect 4154 393932 4160 393984
rect 4212 393972 4218 393984
rect 210694 393972 210700 393984
rect 4212 393944 210700 393972
rect 4212 393932 4218 393944
rect 210694 393932 210700 393944
rect 210752 393932 210758 393984
rect 212626 393932 212632 393984
rect 212684 393972 212690 393984
rect 213178 393972 213184 393984
rect 212684 393944 213184 393972
rect 212684 393932 212690 393944
rect 213178 393932 213184 393944
rect 213236 393932 213242 393984
rect 214006 393932 214012 393984
rect 214064 393972 214070 393984
rect 214834 393972 214840 393984
rect 214064 393944 214840 393972
rect 214064 393932 214070 393944
rect 214834 393932 214840 393944
rect 214892 393932 214898 393984
rect 215662 393932 215668 393984
rect 215720 393972 215726 393984
rect 216030 393972 216036 393984
rect 215720 393944 216036 393972
rect 215720 393932 215726 393944
rect 216030 393932 216036 393944
rect 216088 393932 216094 393984
rect 216858 393932 216864 393984
rect 216916 393972 216922 393984
rect 217594 393972 217600 393984
rect 216916 393944 217600 393972
rect 216916 393932 216922 393944
rect 217594 393932 217600 393944
rect 217652 393932 217658 393984
rect 218606 393932 218612 393984
rect 218664 393972 218670 393984
rect 219066 393972 219072 393984
rect 218664 393944 219072 393972
rect 218664 393932 218670 393944
rect 219066 393932 219072 393944
rect 219124 393932 219130 393984
rect 219802 393932 219808 393984
rect 219860 393972 219866 393984
rect 220262 393972 220268 393984
rect 219860 393944 220268 393972
rect 219860 393932 219866 393944
rect 220262 393932 220268 393944
rect 220320 393932 220326 393984
rect 221090 393932 221096 393984
rect 221148 393972 221154 393984
rect 222102 393972 222108 393984
rect 221148 393944 222108 393972
rect 221148 393932 221154 393944
rect 222102 393932 222108 393944
rect 222160 393932 222166 393984
rect 222470 393932 222476 393984
rect 222528 393972 222534 393984
rect 222930 393972 222936 393984
rect 222528 393944 222936 393972
rect 222528 393932 222534 393944
rect 222930 393932 222936 393944
rect 222988 393932 222994 393984
rect 223850 393932 223856 393984
rect 223908 393972 223914 393984
rect 224862 393972 224868 393984
rect 223908 393944 224868 393972
rect 223908 393932 223914 393944
rect 224862 393932 224868 393944
rect 224920 393932 224926 393984
rect 234982 393932 234988 393984
rect 235040 393972 235046 393984
rect 235350 393972 235356 393984
rect 235040 393944 235356 393972
rect 235040 393932 235046 393944
rect 235350 393932 235356 393944
rect 235408 393932 235414 393984
rect 235994 393932 236000 393984
rect 236052 393972 236058 393984
rect 236638 393972 236644 393984
rect 236052 393944 236644 393972
rect 236052 393932 236058 393944
rect 236638 393932 236644 393944
rect 236696 393932 236702 393984
rect 237576 393916 237604 394216
rect 237742 394204 237748 394216
rect 237800 394204 237806 394256
rect 237852 394244 237880 394352
rect 239508 394244 239536 394352
rect 240134 394272 240140 394324
rect 240192 394312 240198 394324
rect 241440 394312 241468 394352
rect 243998 394340 244004 394392
rect 244056 394380 244062 394392
rect 329834 394380 329840 394392
rect 244056 394352 329840 394380
rect 244056 394340 244062 394352
rect 329834 394340 329840 394352
rect 329892 394340 329898 394392
rect 332594 394312 332600 394324
rect 240192 394284 241376 394312
rect 241440 394284 332600 394312
rect 240192 394272 240198 394284
rect 237852 394216 239536 394244
rect 238846 394136 238852 394188
rect 238904 394176 238910 394188
rect 239398 394176 239404 394188
rect 238904 394148 239404 394176
rect 238904 394136 238910 394148
rect 239398 394136 239404 394148
rect 239456 394136 239462 394188
rect 240134 394136 240140 394188
rect 240192 394176 240198 394188
rect 240686 394176 240692 394188
rect 240192 394148 240692 394176
rect 240192 394136 240198 394148
rect 240686 394136 240692 394148
rect 240744 394136 240750 394188
rect 240226 394068 240232 394120
rect 240284 394108 240290 394120
rect 240594 394108 240600 394120
rect 240284 394080 240600 394108
rect 240284 394068 240290 394080
rect 240594 394068 240600 394080
rect 240652 394068 240658 394120
rect 240318 394000 240324 394052
rect 240376 394040 240382 394052
rect 240686 394040 240692 394052
rect 240376 394012 240692 394040
rect 240376 394000 240382 394012
rect 240686 394000 240692 394012
rect 240744 394000 240750 394052
rect 241348 394040 241376 394284
rect 332594 394272 332600 394284
rect 332652 394272 332658 394324
rect 243170 394204 243176 394256
rect 243228 394244 243234 394256
rect 243538 394244 243544 394256
rect 243228 394216 243544 394244
rect 243228 394204 243234 394216
rect 243538 394204 243544 394216
rect 243596 394204 243602 394256
rect 243906 394204 243912 394256
rect 243964 394244 243970 394256
rect 347774 394244 347780 394256
rect 243964 394216 347780 394244
rect 243964 394204 243970 394216
rect 347774 394204 347780 394216
rect 347832 394204 347838 394256
rect 243354 394136 243360 394188
rect 243412 394176 243418 394188
rect 243722 394176 243728 394188
rect 243412 394148 243728 394176
rect 243412 394136 243418 394148
rect 243722 394136 243728 394148
rect 243780 394136 243786 394188
rect 244366 394136 244372 394188
rect 244424 394176 244430 394188
rect 245194 394176 245200 394188
rect 244424 394148 245200 394176
rect 244424 394136 244430 394148
rect 245194 394136 245200 394148
rect 245252 394136 245258 394188
rect 246206 394136 246212 394188
rect 246264 394176 246270 394188
rect 340874 394176 340880 394188
rect 246264 394148 340880 394176
rect 246264 394136 246270 394148
rect 340874 394136 340880 394148
rect 340932 394136 340938 394188
rect 241514 394068 241520 394120
rect 241572 394108 241578 394120
rect 241882 394108 241888 394120
rect 241572 394080 241888 394108
rect 241572 394068 241578 394080
rect 241882 394068 241888 394080
rect 241940 394068 241946 394120
rect 244274 394068 244280 394120
rect 244332 394108 244338 394120
rect 244918 394108 244924 394120
rect 244332 394080 244924 394108
rect 244332 394068 244338 394080
rect 244918 394068 244924 394080
rect 244976 394068 244982 394120
rect 246942 394068 246948 394120
rect 247000 394108 247006 394120
rect 372614 394108 372620 394120
rect 247000 394080 372620 394108
rect 247000 394068 247006 394080
rect 372614 394068 372620 394080
rect 372672 394068 372678 394120
rect 241348 394012 244596 394040
rect 240594 393932 240600 393984
rect 240652 393972 240658 393984
rect 241054 393972 241060 393984
rect 240652 393944 241060 393972
rect 240652 393932 240658 393944
rect 241054 393932 241060 393944
rect 241112 393932 241118 393984
rect 241606 393932 241612 393984
rect 241664 393972 241670 393984
rect 242158 393972 242164 393984
rect 241664 393944 242164 393972
rect 241664 393932 241670 393944
rect 242158 393932 242164 393944
rect 242216 393932 242222 393984
rect 210142 393864 210148 393916
rect 210200 393904 210206 393916
rect 210602 393904 210608 393916
rect 210200 393876 210608 393904
rect 210200 393864 210206 393876
rect 210602 393864 210608 393876
rect 210660 393864 210666 393916
rect 211430 393864 211436 393916
rect 211488 393904 211494 393916
rect 212074 393904 212080 393916
rect 211488 393876 212080 393904
rect 211488 393864 211494 393876
rect 212074 393864 212080 393876
rect 212132 393864 212138 393916
rect 212810 393864 212816 393916
rect 212868 393904 212874 393916
rect 213822 393904 213828 393916
rect 212868 393876 213828 393904
rect 212868 393864 212874 393876
rect 213822 393864 213828 393876
rect 213880 393864 213886 393916
rect 214558 393864 214564 393916
rect 214616 393904 214622 393916
rect 215202 393904 215208 393916
rect 214616 393876 215208 393904
rect 214616 393864 214622 393876
rect 215202 393864 215208 393876
rect 215260 393864 215266 393916
rect 215478 393864 215484 393916
rect 215536 393904 215542 393916
rect 216214 393904 216220 393916
rect 215536 393876 216220 393904
rect 215536 393864 215542 393876
rect 216214 393864 216220 393876
rect 216272 393864 216278 393916
rect 216766 393864 216772 393916
rect 216824 393904 216830 393916
rect 217870 393904 217876 393916
rect 216824 393876 217876 393904
rect 216824 393864 216830 393876
rect 217870 393864 217876 393876
rect 217928 393864 217934 393916
rect 218330 393864 218336 393916
rect 218388 393904 218394 393916
rect 219250 393904 219256 393916
rect 218388 393876 219256 393904
rect 218388 393864 218394 393876
rect 219250 393864 219256 393876
rect 219308 393864 219314 393916
rect 219710 393864 219716 393916
rect 219768 393904 219774 393916
rect 220630 393904 220636 393916
rect 219768 393876 220636 393904
rect 219768 393864 219774 393876
rect 220630 393864 220636 393876
rect 220688 393864 220694 393916
rect 222746 393864 222752 393916
rect 222804 393904 222810 393916
rect 223206 393904 223212 393916
rect 222804 393876 223212 393904
rect 222804 393864 222810 393876
rect 223206 393864 223212 393876
rect 223264 393864 223270 393916
rect 236178 393864 236184 393916
rect 236236 393904 236242 393916
rect 236236 393876 236316 393904
rect 236236 393864 236242 393876
rect 209958 393796 209964 393848
rect 210016 393836 210022 393848
rect 210510 393836 210516 393848
rect 210016 393808 210516 393836
rect 210016 393796 210022 393808
rect 210510 393796 210516 393808
rect 210568 393796 210574 393848
rect 211614 393796 211620 393848
rect 211672 393836 211678 393848
rect 212350 393836 212356 393848
rect 211672 393808 212356 393836
rect 211672 393796 211678 393808
rect 212350 393796 212356 393808
rect 212408 393796 212414 393848
rect 214374 393796 214380 393848
rect 214432 393836 214438 393848
rect 214926 393836 214932 393848
rect 214432 393808 214932 393836
rect 214432 393796 214438 393808
rect 214926 393796 214932 393808
rect 214984 393796 214990 393848
rect 218514 393796 218520 393848
rect 218572 393836 218578 393848
rect 219158 393836 219164 393848
rect 218572 393808 219164 393836
rect 218572 393796 218578 393808
rect 219158 393796 219164 393808
rect 219216 393796 219222 393848
rect 219894 393796 219900 393848
rect 219952 393836 219958 393848
rect 220722 393836 220728 393848
rect 219952 393808 220728 393836
rect 219952 393796 219958 393808
rect 220722 393796 220728 393808
rect 220780 393796 220786 393848
rect 224034 393796 224040 393848
rect 224092 393836 224098 393848
rect 224310 393836 224316 393848
rect 224092 393808 224316 393836
rect 224092 393796 224098 393808
rect 224310 393796 224316 393808
rect 224368 393796 224374 393848
rect 234798 393796 234804 393848
rect 234856 393836 234862 393848
rect 235718 393836 235724 393848
rect 234856 393808 235724 393836
rect 234856 393796 234862 393808
rect 235718 393796 235724 393808
rect 235776 393796 235782 393848
rect 214098 393728 214104 393780
rect 214156 393768 214162 393780
rect 215110 393768 215116 393780
rect 214156 393740 215116 393768
rect 214156 393728 214162 393740
rect 215110 393728 215116 393740
rect 215168 393728 215174 393780
rect 221182 393728 221188 393780
rect 221240 393768 221246 393780
rect 221826 393768 221832 393780
rect 221240 393740 221832 393768
rect 221240 393728 221246 393740
rect 221826 393728 221832 393740
rect 221884 393728 221890 393780
rect 236288 393712 236316 393876
rect 237558 393864 237564 393916
rect 237616 393864 237622 393916
rect 240410 393864 240416 393916
rect 240468 393904 240474 393916
rect 241238 393904 241244 393916
rect 240468 393876 241244 393904
rect 240468 393864 240474 393876
rect 241238 393864 241244 393876
rect 241296 393864 241302 393916
rect 241882 393864 241888 393916
rect 241940 393904 241946 393916
rect 242342 393904 242348 393916
rect 241940 393876 242348 393904
rect 241940 393864 241946 393876
rect 242342 393864 242348 393876
rect 242400 393864 242406 393916
rect 243078 393864 243084 393916
rect 243136 393904 243142 393916
rect 243446 393904 243452 393916
rect 243136 393876 243452 393904
rect 243136 393864 243142 393876
rect 243446 393864 243452 393876
rect 243504 393864 243510 393916
rect 244568 393904 244596 394012
rect 244642 394000 244648 394052
rect 244700 394040 244706 394052
rect 245194 394040 245200 394052
rect 244700 394012 245200 394040
rect 244700 394000 244706 394012
rect 245194 394000 245200 394012
rect 245252 394000 245258 394052
rect 249886 394000 249892 394052
rect 249944 394040 249950 394052
rect 250530 394040 250536 394052
rect 249944 394012 250536 394040
rect 249944 394000 249950 394012
rect 250530 394000 250536 394012
rect 250588 394000 250594 394052
rect 252830 394000 252836 394052
rect 252888 394040 252894 394052
rect 253198 394040 253204 394052
rect 252888 394012 253204 394040
rect 252888 394000 252894 394012
rect 253198 394000 253204 394012
rect 253256 394000 253262 394052
rect 382274 394040 382280 394052
rect 253906 394012 382280 394040
rect 251542 393932 251548 393984
rect 251600 393972 251606 393984
rect 251726 393972 251732 393984
rect 251600 393944 251732 393972
rect 251600 393932 251606 393944
rect 251726 393932 251732 393944
rect 251784 393932 251790 393984
rect 252646 393932 252652 393984
rect 252704 393972 252710 393984
rect 252922 393972 252928 393984
rect 252704 393944 252928 393972
rect 252704 393932 252710 393944
rect 252922 393932 252928 393944
rect 252980 393932 252986 393984
rect 253906 393904 253934 394012
rect 382274 394000 382280 394012
rect 382332 394000 382338 394052
rect 254762 393932 254768 393984
rect 254820 393972 254826 393984
rect 571334 393972 571340 393984
rect 254820 393944 571340 393972
rect 254820 393932 254826 393944
rect 571334 393932 571340 393944
rect 571392 393932 571398 393984
rect 244568 393876 253934 393904
rect 237374 393796 237380 393848
rect 237432 393836 237438 393848
rect 238294 393836 238300 393848
rect 237432 393808 238300 393836
rect 237432 393796 237438 393808
rect 238294 393796 238300 393808
rect 238352 393796 238358 393848
rect 240318 393796 240324 393848
rect 240376 393836 240382 393848
rect 241146 393836 241152 393848
rect 240376 393808 241152 393836
rect 240376 393796 240382 393808
rect 241146 393796 241152 393808
rect 241204 393796 241210 393848
rect 241698 393796 241704 393848
rect 241756 393836 241762 393848
rect 241974 393836 241980 393848
rect 241756 393808 241980 393836
rect 241756 393796 241762 393808
rect 241974 393796 241980 393808
rect 242032 393796 242038 393848
rect 244458 393796 244464 393848
rect 244516 393836 244522 393848
rect 244734 393836 244740 393848
rect 244516 393808 244740 393836
rect 244516 393796 244522 393808
rect 244734 393796 244740 393808
rect 244792 393796 244798 393848
rect 247034 393796 247040 393848
rect 247092 393836 247098 393848
rect 247310 393836 247316 393848
rect 247092 393808 247316 393836
rect 247092 393796 247098 393808
rect 247310 393796 247316 393808
rect 247368 393796 247374 393848
rect 247402 393796 247408 393848
rect 247460 393836 247466 393848
rect 247862 393836 247868 393848
rect 247460 393808 247868 393836
rect 247460 393796 247466 393808
rect 247862 393796 247868 393808
rect 247920 393796 247926 393848
rect 248690 393796 248696 393848
rect 248748 393836 248754 393848
rect 248966 393836 248972 393848
rect 248748 393808 248972 393836
rect 248748 393796 248754 393808
rect 248966 393796 248972 393808
rect 249024 393796 249030 393848
rect 249978 393796 249984 393848
rect 250036 393836 250042 393848
rect 250254 393836 250260 393848
rect 250036 393808 250260 393836
rect 250036 393796 250042 393808
rect 250254 393796 250260 393808
rect 250312 393796 250318 393848
rect 251174 393796 251180 393848
rect 251232 393836 251238 393848
rect 251726 393836 251732 393848
rect 251232 393808 251732 393836
rect 251232 393796 251238 393808
rect 251726 393796 251732 393808
rect 251784 393796 251790 393848
rect 252922 393796 252928 393848
rect 252980 393836 252986 393848
rect 253290 393836 253296 393848
rect 252980 393808 253296 393836
rect 252980 393796 252986 393808
rect 253290 393796 253296 393808
rect 253348 393796 253354 393848
rect 236822 393728 236828 393780
rect 236880 393768 236886 393780
rect 244182 393768 244188 393780
rect 236880 393740 244188 393768
rect 236880 393728 236886 393740
rect 244182 393728 244188 393740
rect 244240 393728 244246 393780
rect 244550 393728 244556 393780
rect 244608 393768 244614 393780
rect 245286 393768 245292 393780
rect 244608 393740 245292 393768
rect 244608 393728 244614 393740
rect 245286 393728 245292 393740
rect 245344 393728 245350 393780
rect 252830 393728 252836 393780
rect 252888 393768 252894 393780
rect 253382 393768 253388 393780
rect 252888 393740 253388 393768
rect 252888 393728 252894 393740
rect 253382 393728 253388 393740
rect 253440 393728 253446 393780
rect 213086 393660 213092 393712
rect 213144 393700 213150 393712
rect 213638 393700 213644 393712
rect 213144 393672 213644 393700
rect 213144 393660 213150 393672
rect 213638 393660 213644 393672
rect 213696 393660 213702 393712
rect 235258 393660 235264 393712
rect 235316 393700 235322 393712
rect 235442 393700 235448 393712
rect 235316 393672 235448 393700
rect 235316 393660 235322 393672
rect 235442 393660 235448 393672
rect 235500 393660 235506 393712
rect 236270 393660 236276 393712
rect 236328 393660 236334 393712
rect 236362 393660 236368 393712
rect 236420 393700 236426 393712
rect 236914 393700 236920 393712
rect 236420 393672 236920 393700
rect 236420 393660 236426 393672
rect 236914 393660 236920 393672
rect 236972 393660 236978 393712
rect 243170 393660 243176 393712
rect 243228 393700 243234 393712
rect 243814 393700 243820 393712
rect 243228 393672 243820 393700
rect 243228 393660 243234 393672
rect 243814 393660 243820 393672
rect 243872 393660 243878 393712
rect 244734 393660 244740 393712
rect 244792 393700 244798 393712
rect 245010 393700 245016 393712
rect 244792 393672 245016 393700
rect 244792 393660 244798 393672
rect 245010 393660 245016 393672
rect 245068 393660 245074 393712
rect 251174 393660 251180 393712
rect 251232 393700 251238 393712
rect 251818 393700 251824 393712
rect 251232 393672 251824 393700
rect 251232 393660 251238 393672
rect 251818 393660 251824 393672
rect 251876 393660 251882 393712
rect 244826 393592 244832 393644
rect 244884 393632 244890 393644
rect 244884 393604 244964 393632
rect 244884 393592 244890 393604
rect 244936 393440 244964 393604
rect 244918 393388 244924 393440
rect 244976 393388 244982 393440
rect 227898 393320 227904 393372
rect 227956 393360 227962 393372
rect 228450 393360 228456 393372
rect 227956 393332 228456 393360
rect 227956 393320 227962 393332
rect 228450 393320 228456 393332
rect 228508 393320 228514 393372
rect 221458 393184 221464 393236
rect 221516 393224 221522 393236
rect 221918 393224 221924 393236
rect 221516 393196 221924 393224
rect 221516 393184 221522 393196
rect 221918 393184 221924 393196
rect 221976 393184 221982 393236
rect 239858 392776 239864 392828
rect 239916 392816 239922 392828
rect 277394 392816 277400 392828
rect 239916 392788 277400 392816
rect 239916 392776 239922 392788
rect 277394 392776 277400 392788
rect 277452 392776 277458 392828
rect 232590 392708 232596 392760
rect 232648 392748 232654 392760
rect 281534 392748 281540 392760
rect 232648 392720 281540 392748
rect 232648 392708 232654 392720
rect 281534 392708 281540 392720
rect 281592 392708 281598 392760
rect 160094 392640 160100 392692
rect 160152 392680 160158 392692
rect 217778 392680 217784 392692
rect 160152 392652 217784 392680
rect 160152 392640 160158 392652
rect 217778 392640 217784 392652
rect 217836 392640 217842 392692
rect 242434 392640 242440 392692
rect 242492 392680 242498 392692
rect 401594 392680 401600 392692
rect 242492 392652 401600 392680
rect 242492 392640 242498 392652
rect 401594 392640 401600 392652
rect 401652 392640 401658 392692
rect 109034 392572 109040 392624
rect 109092 392612 109098 392624
rect 218882 392612 218888 392624
rect 109092 392584 218888 392612
rect 109092 392572 109098 392584
rect 218882 392572 218888 392584
rect 218940 392572 218946 392624
rect 249242 392572 249248 392624
rect 249300 392612 249306 392624
rect 498194 392612 498200 392624
rect 249300 392584 498200 392612
rect 249300 392572 249306 392584
rect 498194 392572 498200 392584
rect 498252 392572 498258 392624
rect 218698 392504 218704 392556
rect 218756 392544 218762 392556
rect 218756 392516 218836 392544
rect 218756 392504 218762 392516
rect 218808 392352 218836 392516
rect 245654 392368 245660 392420
rect 245712 392408 245718 392420
rect 246206 392408 246212 392420
rect 245712 392380 246212 392408
rect 245712 392368 245718 392380
rect 246206 392368 246212 392380
rect 246264 392368 246270 392420
rect 218790 392300 218796 392352
rect 218848 392300 218854 392352
rect 210050 392164 210056 392216
rect 210108 392204 210114 392216
rect 210878 392204 210884 392216
rect 210108 392176 210884 392204
rect 210108 392164 210114 392176
rect 210878 392164 210884 392176
rect 210936 392164 210942 392216
rect 222930 392164 222936 392216
rect 222988 392204 222994 392216
rect 223298 392204 223304 392216
rect 222988 392176 223304 392204
rect 222988 392164 222994 392176
rect 223298 392164 223304 392176
rect 223356 392164 223362 392216
rect 245746 392164 245752 392216
rect 245804 392204 245810 392216
rect 246298 392204 246304 392216
rect 245804 392176 246304 392204
rect 245804 392164 245810 392176
rect 246298 392164 246304 392176
rect 246356 392164 246362 392216
rect 238938 392096 238944 392148
rect 238996 392136 239002 392148
rect 239674 392136 239680 392148
rect 238996 392108 239680 392136
rect 238996 392096 239002 392108
rect 239674 392096 239680 392108
rect 239732 392096 239738 392148
rect 250254 392096 250260 392148
rect 250312 392136 250318 392148
rect 250438 392136 250444 392148
rect 250312 392108 250444 392136
rect 250312 392096 250318 392108
rect 250438 392096 250444 392108
rect 250496 392096 250502 392148
rect 247126 392028 247132 392080
rect 247184 392068 247190 392080
rect 247770 392068 247776 392080
rect 247184 392040 247776 392068
rect 247184 392028 247190 392040
rect 247770 392028 247776 392040
rect 247828 392028 247834 392080
rect 248414 392028 248420 392080
rect 248472 392068 248478 392080
rect 248874 392068 248880 392080
rect 248472 392040 248880 392068
rect 248472 392028 248478 392040
rect 248874 392028 248880 392040
rect 248932 392028 248938 392080
rect 249794 392028 249800 392080
rect 249852 392068 249858 392080
rect 250162 392068 250168 392080
rect 249852 392040 250168 392068
rect 249852 392028 249858 392040
rect 250162 392028 250168 392040
rect 250220 392028 250226 392080
rect 248690 391960 248696 392012
rect 248748 392000 248754 392012
rect 249426 392000 249432 392012
rect 248748 391972 249432 392000
rect 248748 391960 248754 391972
rect 249426 391960 249432 391972
rect 249484 391960 249490 392012
rect 248414 391892 248420 391944
rect 248472 391932 248478 391944
rect 249334 391932 249340 391944
rect 248472 391904 249340 391932
rect 248472 391892 248478 391904
rect 249334 391892 249340 391904
rect 249392 391892 249398 391944
rect 249794 391892 249800 391944
rect 249852 391932 249858 391944
rect 250714 391932 250720 391944
rect 249852 391904 250720 391932
rect 249852 391892 249858 391904
rect 250714 391892 250720 391904
rect 250772 391892 250778 391944
rect 216398 391864 216404 391876
rect 216048 391836 216404 391864
rect 216048 391808 216076 391836
rect 216398 391824 216404 391836
rect 216456 391824 216462 391876
rect 216030 391756 216036 391808
rect 216088 391756 216094 391808
rect 215846 391620 215852 391672
rect 215904 391660 215910 391672
rect 216214 391660 216220 391672
rect 215904 391632 216220 391660
rect 215904 391620 215910 391632
rect 216214 391620 216220 391632
rect 216272 391620 216278 391672
rect 238202 391552 238208 391604
rect 238260 391592 238266 391604
rect 331214 391592 331220 391604
rect 238260 391564 331220 391592
rect 238260 391552 238266 391564
rect 331214 391552 331220 391564
rect 331272 391552 331278 391604
rect 215846 391484 215852 391536
rect 215904 391524 215910 391536
rect 216582 391524 216588 391536
rect 215904 391496 216588 391524
rect 215904 391484 215910 391496
rect 216582 391484 216588 391496
rect 216640 391484 216646 391536
rect 239766 391484 239772 391536
rect 239824 391524 239830 391536
rect 365714 391524 365720 391536
rect 239824 391496 365720 391524
rect 239824 391484 239830 391496
rect 365714 391484 365720 391496
rect 365772 391484 365778 391536
rect 247954 391416 247960 391468
rect 248012 391456 248018 391468
rect 387794 391456 387800 391468
rect 248012 391428 387800 391456
rect 248012 391416 248018 391428
rect 387794 391416 387800 391428
rect 387852 391416 387858 391468
rect 245378 391348 245384 391400
rect 245436 391388 245442 391400
rect 440234 391388 440240 391400
rect 245436 391360 440240 391388
rect 245436 391348 245442 391360
rect 440234 391348 440240 391360
rect 440292 391348 440298 391400
rect 245838 391280 245844 391332
rect 245896 391320 245902 391332
rect 456794 391320 456800 391332
rect 245896 391292 456800 391320
rect 245896 391280 245902 391292
rect 456794 391280 456800 391292
rect 456852 391280 456858 391332
rect 210326 391212 210332 391264
rect 210384 391252 210390 391264
rect 210510 391252 210516 391264
rect 210384 391224 210516 391252
rect 210384 391212 210390 391224
rect 210510 391212 210516 391224
rect 210568 391212 210574 391264
rect 237834 391212 237840 391264
rect 237892 391252 237898 391264
rect 238386 391252 238392 391264
rect 237892 391224 238392 391252
rect 237892 391212 237898 391224
rect 238386 391212 238392 391224
rect 238444 391212 238450 391264
rect 250806 391212 250812 391264
rect 250864 391252 250870 391264
rect 511994 391252 512000 391264
rect 250864 391224 512000 391252
rect 250864 391212 250870 391224
rect 511994 391212 512000 391224
rect 512052 391212 512058 391264
rect 245838 391008 245844 391060
rect 245896 391048 245902 391060
rect 246574 391048 246580 391060
rect 245896 391020 246580 391048
rect 245896 391008 245902 391020
rect 246574 391008 246580 391020
rect 246632 391008 246638 391060
rect 239214 390600 239220 390652
rect 239272 390640 239278 390652
rect 239490 390640 239496 390652
rect 239272 390612 239496 390640
rect 239272 390600 239278 390612
rect 239490 390600 239496 390612
rect 239548 390600 239554 390652
rect 210234 390532 210240 390584
rect 210292 390572 210298 390584
rect 210970 390572 210976 390584
rect 210292 390544 210976 390572
rect 210292 390532 210298 390544
rect 210970 390532 210976 390544
rect 211028 390532 211034 390584
rect 210326 390464 210332 390516
rect 210384 390504 210390 390516
rect 211062 390504 211068 390516
rect 210384 390476 211068 390504
rect 210384 390464 210390 390476
rect 211062 390464 211068 390476
rect 211120 390464 211126 390516
rect 251266 390464 251272 390516
rect 251324 390504 251330 390516
rect 252094 390504 252100 390516
rect 251324 390476 252100 390504
rect 251324 390464 251330 390476
rect 252094 390464 252100 390476
rect 252152 390464 252158 390516
rect 214466 390396 214472 390448
rect 214524 390436 214530 390448
rect 214742 390436 214748 390448
rect 214524 390408 214748 390436
rect 214524 390396 214530 390408
rect 214742 390396 214748 390408
rect 214800 390396 214806 390448
rect 217226 390260 217232 390312
rect 217284 390300 217290 390312
rect 217502 390300 217508 390312
rect 217284 390272 217508 390300
rect 217284 390260 217290 390272
rect 217502 390260 217508 390272
rect 217560 390260 217566 390312
rect 246114 390056 246120 390108
rect 246172 390096 246178 390108
rect 246390 390096 246396 390108
rect 246172 390068 246396 390096
rect 246172 390056 246178 390068
rect 246390 390056 246396 390068
rect 246448 390056 246454 390108
rect 222562 389988 222568 390040
rect 222620 390028 222626 390040
rect 223206 390028 223212 390040
rect 222620 390000 223212 390028
rect 222620 389988 222626 390000
rect 223206 389988 223212 390000
rect 223264 389988 223270 390040
rect 233970 389920 233976 389972
rect 234028 389960 234034 389972
rect 298094 389960 298100 389972
rect 234028 389932 298100 389960
rect 234028 389920 234034 389932
rect 298094 389920 298100 389932
rect 298152 389920 298158 389972
rect 222562 389852 222568 389904
rect 222620 389892 222626 389904
rect 223482 389892 223488 389904
rect 222620 389864 223488 389892
rect 222620 389852 222626 389864
rect 223482 389852 223488 389864
rect 223540 389852 223546 389904
rect 240870 389852 240876 389904
rect 240928 389892 240934 389904
rect 391934 389892 391940 389904
rect 240928 389864 391940 389892
rect 240928 389852 240934 389864
rect 391934 389852 391940 389864
rect 391992 389852 391998 389904
rect 223758 389784 223764 389836
rect 223816 389824 223822 389836
rect 224586 389824 224592 389836
rect 223816 389796 224592 389824
rect 223816 389784 223822 389796
rect 224586 389784 224592 389796
rect 224644 389784 224650 389836
rect 249518 389784 249524 389836
rect 249576 389824 249582 389836
rect 499574 389824 499580 389836
rect 249576 389796 499580 389824
rect 249576 389784 249582 389796
rect 499574 389784 499580 389796
rect 499632 389784 499638 389836
rect 250438 389308 250444 389360
rect 250496 389348 250502 389360
rect 250622 389348 250628 389360
rect 250496 389320 250628 389348
rect 250496 389308 250502 389320
rect 250622 389308 250628 389320
rect 250680 389308 250686 389360
rect 299198 379448 299204 379500
rect 299256 379488 299262 379500
rect 580166 379488 580172 379500
rect 299256 379460 580172 379488
rect 299256 379448 299262 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 98638 372552 98644 372564
rect 3384 372524 98644 372552
rect 3384 372512 3390 372524
rect 98638 372512 98644 372524
rect 98696 372512 98702 372564
rect 295886 365644 295892 365696
rect 295944 365684 295950 365696
rect 580166 365684 580172 365696
rect 295944 365656 580172 365684
rect 295944 365644 295950 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 106274 363604 106280 363656
rect 106332 363644 106338 363656
rect 209314 363644 209320 363656
rect 106332 363616 209320 363644
rect 106332 363604 106338 363616
rect 209314 363604 209320 363616
rect 209372 363604 209378 363656
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4890 358476 4896 358488
rect 2832 358448 4896 358476
rect 2832 358436 2838 358448
rect 4890 358436 4896 358448
rect 4948 358436 4954 358488
rect 92474 355444 92480 355496
rect 92532 355484 92538 355496
rect 217226 355484 217232 355496
rect 92532 355456 217232 355484
rect 92532 355444 92538 355456
rect 217226 355444 217232 355456
rect 217284 355444 217290 355496
rect 232498 355444 232504 355496
rect 232556 355484 232562 355496
rect 284294 355484 284300 355496
rect 232556 355456 284300 355484
rect 232556 355444 232562 355456
rect 284294 355444 284300 355456
rect 284352 355444 284358 355496
rect 42794 355376 42800 355428
rect 42852 355416 42858 355428
rect 213086 355416 213092 355428
rect 42852 355388 213092 355416
rect 42852 355376 42858 355388
rect 213086 355376 213092 355388
rect 213144 355376 213150 355428
rect 244734 355376 244740 355428
rect 244792 355416 244798 355428
rect 445754 355416 445760 355428
rect 244792 355388 445760 355416
rect 244792 355376 244798 355388
rect 445754 355376 445760 355388
rect 445812 355376 445818 355428
rect 37274 355308 37280 355360
rect 37332 355348 37338 355360
rect 212994 355348 213000 355360
rect 37332 355320 213000 355348
rect 37332 355308 37338 355320
rect 212994 355308 213000 355320
rect 213052 355308 213058 355360
rect 250530 355308 250536 355360
rect 250588 355348 250594 355360
rect 514754 355348 514760 355360
rect 250588 355320 514760 355348
rect 250588 355308 250594 355320
rect 514754 355308 514760 355320
rect 514812 355308 514818 355360
rect 169018 354424 169024 354476
rect 169076 354464 169082 354476
rect 218606 354464 218612 354476
rect 169076 354436 218612 354464
rect 169076 354424 169082 354436
rect 218606 354424 218612 354436
rect 218664 354424 218670 354476
rect 88334 354356 88340 354408
rect 88392 354396 88398 354408
rect 213178 354396 213184 354408
rect 88392 354368 213184 354396
rect 88392 354356 88398 354368
rect 213178 354356 213184 354368
rect 213236 354356 213242 354408
rect 91094 354288 91100 354340
rect 91152 354328 91158 354340
rect 217042 354328 217048 354340
rect 91152 354300 217048 354328
rect 91152 354288 91158 354300
rect 217042 354288 217048 354300
rect 217100 354288 217106 354340
rect 231026 354288 231032 354340
rect 231084 354328 231090 354340
rect 262214 354328 262220 354340
rect 231084 354300 262220 354328
rect 231084 354288 231090 354300
rect 262214 354288 262220 354300
rect 262272 354288 262278 354340
rect 86954 354220 86960 354272
rect 87012 354260 87018 354272
rect 217134 354260 217140 354272
rect 87012 354232 217140 354260
rect 87012 354220 87018 354232
rect 217134 354220 217140 354232
rect 217192 354220 217198 354272
rect 246574 354220 246580 354272
rect 246632 354260 246638 354272
rect 357434 354260 357440 354272
rect 246632 354232 357440 354260
rect 246632 354220 246638 354232
rect 357434 354220 357440 354232
rect 357492 354220 357498 354272
rect 70394 354152 70400 354204
rect 70452 354192 70458 354204
rect 212074 354192 212080 354204
rect 70452 354164 212080 354192
rect 70452 354152 70458 354164
rect 212074 354152 212080 354164
rect 212132 354152 212138 354204
rect 240870 354152 240876 354204
rect 240928 354192 240934 354204
rect 393314 354192 393320 354204
rect 240928 354164 393320 354192
rect 240928 354152 240934 354164
rect 393314 354152 393320 354164
rect 393372 354152 393378 354204
rect 60734 354084 60740 354136
rect 60792 354124 60798 354136
rect 211982 354124 211988 354136
rect 60792 354096 211988 354124
rect 60792 354084 60798 354096
rect 211982 354084 211988 354096
rect 212040 354084 212046 354136
rect 228358 354084 228364 354136
rect 228416 354124 228422 354136
rect 232498 354124 232504 354136
rect 228416 354096 232504 354124
rect 228416 354084 228422 354096
rect 232498 354084 232504 354096
rect 232556 354084 232562 354136
rect 245010 354084 245016 354136
rect 245068 354124 245074 354136
rect 440326 354124 440332 354136
rect 245068 354096 440332 354124
rect 245068 354084 245074 354096
rect 440326 354084 440332 354096
rect 440384 354084 440390 354136
rect 62114 354016 62120 354068
rect 62172 354056 62178 354068
rect 214558 354056 214564 354068
rect 62172 354028 214564 354056
rect 62172 354016 62178 354028
rect 214558 354016 214564 354028
rect 214616 354016 214622 354068
rect 229738 354016 229744 354068
rect 229796 354056 229802 354068
rect 240778 354056 240784 354068
rect 229796 354028 240784 354056
rect 229796 354016 229802 354028
rect 240778 354016 240784 354028
rect 240836 354016 240842 354068
rect 251818 354016 251824 354068
rect 251876 354056 251882 354068
rect 534074 354056 534080 354068
rect 251876 354028 534080 354056
rect 251876 354016 251882 354028
rect 534074 354016 534080 354028
rect 534132 354016 534138 354068
rect 56594 353948 56600 354000
rect 56652 353988 56658 354000
rect 214466 353988 214472 354000
rect 56652 353960 214472 353988
rect 56652 353948 56658 353960
rect 214466 353948 214472 353960
rect 214524 353948 214530 354000
rect 229830 353948 229836 354000
rect 229888 353988 229894 354000
rect 244734 353988 244740 354000
rect 229888 353960 244740 353988
rect 229888 353948 229894 353960
rect 244734 353948 244740 353960
rect 244792 353948 244798 354000
rect 253198 353948 253204 354000
rect 253256 353988 253262 354000
rect 546494 353988 546500 354000
rect 253256 353960 546500 353988
rect 253256 353948 253262 353960
rect 546494 353948 546500 353960
rect 546552 353948 546558 354000
rect 299290 353200 299296 353252
rect 299348 353240 299354 353252
rect 580166 353240 580172 353252
rect 299348 353212 580172 353240
rect 299348 353200 299354 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 198734 352724 198740 352776
rect 198792 352764 198798 352776
rect 225506 352764 225512 352776
rect 198792 352736 225512 352764
rect 198792 352724 198798 352736
rect 225506 352724 225512 352736
rect 225564 352724 225570 352776
rect 180794 352656 180800 352708
rect 180852 352696 180858 352708
rect 224218 352696 224224 352708
rect 180852 352668 224224 352696
rect 180852 352656 180858 352668
rect 224218 352656 224224 352668
rect 224276 352656 224282 352708
rect 235350 352656 235356 352708
rect 235408 352696 235414 352708
rect 316034 352696 316040 352708
rect 235408 352668 316040 352696
rect 235408 352656 235414 352668
rect 316034 352656 316040 352668
rect 316092 352656 316098 352708
rect 160186 352588 160192 352640
rect 160244 352628 160250 352640
rect 223022 352628 223028 352640
rect 160244 352600 223028 352628
rect 160244 352588 160250 352600
rect 223022 352588 223028 352600
rect 223080 352588 223086 352640
rect 240686 352588 240692 352640
rect 240744 352628 240750 352640
rect 385034 352628 385040 352640
rect 240744 352600 385040 352628
rect 240744 352588 240750 352600
rect 385034 352588 385040 352600
rect 385092 352588 385098 352640
rect 5534 352520 5540 352572
rect 5592 352560 5598 352572
rect 210418 352560 210424 352572
rect 5592 352532 210424 352560
rect 5592 352520 5598 352532
rect 210418 352520 210424 352532
rect 210476 352520 210482 352572
rect 243630 352520 243636 352572
rect 243688 352560 243694 352572
rect 423674 352560 423680 352572
rect 243688 352532 423680 352560
rect 243688 352520 243694 352532
rect 423674 352520 423680 352532
rect 423732 352520 423738 352572
rect 225690 351908 225696 351960
rect 225748 351948 225754 351960
rect 226886 351948 226892 351960
rect 225748 351920 226892 351948
rect 225748 351908 225754 351920
rect 226886 351908 226892 351920
rect 226944 351908 226950 351960
rect 238110 351228 238116 351280
rect 238168 351268 238174 351280
rect 357526 351268 357532 351280
rect 238168 351240 357532 351268
rect 238168 351228 238174 351240
rect 357526 351228 357532 351240
rect 357584 351228 357590 351280
rect 85574 351160 85580 351212
rect 85632 351200 85638 351212
rect 210510 351200 210516 351212
rect 85632 351172 210516 351200
rect 85632 351160 85638 351172
rect 210510 351160 210516 351172
rect 210568 351160 210574 351212
rect 254578 351160 254584 351212
rect 254636 351200 254642 351212
rect 572714 351200 572720 351212
rect 254636 351172 572720 351200
rect 254636 351160 254642 351172
rect 572714 351160 572720 351172
rect 572772 351160 572778 351212
rect 110414 340144 110420 340196
rect 110472 340184 110478 340196
rect 208026 340184 208032 340196
rect 110472 340156 208032 340184
rect 110472 340144 110478 340156
rect 208026 340144 208032 340156
rect 208084 340144 208090 340196
rect 23474 338716 23480 338768
rect 23532 338756 23538 338768
rect 209222 338756 209228 338768
rect 23532 338728 209228 338756
rect 23532 338716 23538 338728
rect 209222 338716 209228 338728
rect 209280 338716 209286 338768
rect 258810 334568 258816 334620
rect 258868 334608 258874 334620
rect 580994 334608 581000 334620
rect 258868 334580 581000 334608
rect 258868 334568 258874 334580
rect 580994 334568 581000 334580
rect 581052 334568 581058 334620
rect 24854 333208 24860 333260
rect 24912 333248 24918 333260
rect 209130 333248 209136 333260
rect 24912 333220 209136 333248
rect 24912 333208 24918 333220
rect 209130 333208 209136 333220
rect 209188 333208 209194 333260
rect 258718 333208 258724 333260
rect 258776 333248 258782 333260
rect 436094 333248 436100 333260
rect 258776 333220 436100 333248
rect 258776 333208 258782 333220
rect 436094 333208 436100 333220
rect 436152 333208 436158 333260
rect 296622 325592 296628 325644
rect 296680 325632 296686 325644
rect 580166 325632 580172 325644
rect 296680 325604 580172 325632
rect 296680 325592 296686 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 199562 320124 199568 320136
rect 3384 320096 199568 320124
rect 3384 320084 3390 320096
rect 199562 320084 199568 320096
rect 199620 320084 199626 320136
rect 296530 313216 296536 313268
rect 296588 313256 296594 313268
rect 580166 313256 580172 313268
rect 296588 313228 580172 313256
rect 296588 313216 296594 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 200942 306320 200948 306332
rect 3384 306292 200948 306320
rect 3384 306280 3390 306292
rect 200942 306280 200948 306292
rect 201000 306280 201006 306332
rect 257522 304240 257528 304292
rect 257580 304280 257586 304292
rect 429194 304280 429200 304292
rect 257580 304252 429200 304280
rect 257580 304240 257586 304252
rect 429194 304240 429200 304252
rect 429252 304240 429258 304292
rect 265710 299412 265716 299464
rect 265768 299452 265774 299464
rect 580166 299452 580172 299464
rect 265768 299424 580172 299452
rect 265768 299412 265774 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 296438 273164 296444 273216
rect 296496 273204 296502 273216
rect 580166 273204 580172 273216
rect 296496 273176 580172 273204
rect 296496 273164 296502 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3142 267656 3148 267708
rect 3200 267696 3206 267708
rect 196710 267696 196716 267708
rect 3200 267668 196716 267696
rect 3200 267656 3206 267668
rect 196710 267656 196716 267668
rect 196768 267656 196774 267708
rect 296346 259360 296352 259412
rect 296404 259400 296410 259412
rect 580166 259400 580172 259412
rect 296404 259372 580172 259400
rect 296404 259360 296410 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 299106 245556 299112 245608
rect 299164 245596 299170 245608
rect 580166 245596 580172 245608
rect 299164 245568 580172 245596
rect 299164 245556 299170 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 299014 233180 299020 233232
rect 299072 233220 299078 233232
rect 579982 233220 579988 233232
rect 299072 233192 579988 233220
rect 299072 233180 299078 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 296254 219376 296260 219428
rect 296312 219416 296318 219428
rect 580166 219416 580172 219428
rect 296312 219388 580172 219416
rect 296312 219376 296318 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3050 215228 3056 215280
rect 3108 215268 3114 215280
rect 199470 215268 199476 215280
rect 3108 215240 199476 215268
rect 3108 215228 3114 215240
rect 199470 215228 199476 215240
rect 199528 215228 199534 215280
rect 269850 206932 269856 206984
rect 269908 206972 269914 206984
rect 579798 206972 579804 206984
rect 269908 206944 579804 206972
rect 269908 206932 269914 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 271230 193128 271236 193180
rect 271288 193168 271294 193180
rect 580166 193168 580172 193180
rect 271288 193140 580172 193168
rect 271288 193128 271294 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 275278 185580 275284 185632
rect 275336 185620 275342 185632
rect 582374 185620 582380 185632
rect 275336 185592 582380 185620
rect 275336 185580 275342 185592
rect 582374 185580 582380 185592
rect 582432 185580 582438 185632
rect 274082 184152 274088 184204
rect 274140 184192 274146 184204
rect 474734 184192 474740 184204
rect 274140 184164 474740 184192
rect 274140 184152 274146 184164
rect 474734 184152 474740 184164
rect 474792 184152 474798 184204
rect 264330 182792 264336 182844
rect 264388 182832 264394 182844
rect 449894 182832 449900 182844
rect 264388 182804 449900 182832
rect 264388 182792 264394 182804
rect 449894 182792 449900 182804
rect 449952 182792 449958 182844
rect 38654 181432 38660 181484
rect 38712 181472 38718 181484
rect 202138 181472 202144 181484
rect 38712 181444 202144 181472
rect 38712 181432 38718 181444
rect 202138 181432 202144 181444
rect 202196 181432 202202 181484
rect 102226 180072 102232 180124
rect 102284 180112 102290 180124
rect 207934 180112 207940 180124
rect 102284 180084 207940 180112
rect 102284 180072 102290 180084
rect 207934 180072 207940 180084
rect 207992 180072 207998 180124
rect 261478 180072 261484 180124
rect 261536 180112 261542 180124
rect 442994 180112 443000 180124
rect 261536 180084 443000 180112
rect 261536 180072 261542 180084
rect 442994 180072 443000 180084
rect 443052 180072 443058 180124
rect 296162 179324 296168 179376
rect 296220 179364 296226 179376
rect 580166 179364 580172 179376
rect 296220 179336 580172 179364
rect 296220 179324 296226 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 176654 178712 176660 178764
rect 176712 178752 176718 178764
rect 224126 178752 224132 178764
rect 176712 178724 224132 178752
rect 176712 178712 176718 178724
rect 224126 178712 224132 178724
rect 224184 178712 224190 178764
rect 41414 178644 41420 178696
rect 41472 178684 41478 178696
rect 211890 178684 211896 178696
rect 41472 178656 211896 178684
rect 41472 178644 41478 178656
rect 211890 178644 211896 178656
rect 211948 178644 211954 178696
rect 166994 177556 167000 177608
rect 167052 177596 167058 177608
rect 222930 177596 222936 177608
rect 167052 177568 222936 177596
rect 167052 177556 167058 177568
rect 222930 177556 222936 177568
rect 222988 177556 222994 177608
rect 154574 177488 154580 177540
rect 154632 177528 154638 177540
rect 216030 177528 216036 177540
rect 154632 177500 216036 177528
rect 154632 177488 154638 177500
rect 216030 177488 216036 177500
rect 216088 177488 216094 177540
rect 217042 177488 217048 177540
rect 217100 177528 217106 177540
rect 226702 177528 226708 177540
rect 217100 177500 226708 177528
rect 217100 177488 217106 177500
rect 226702 177488 226708 177500
rect 226760 177488 226766 177540
rect 140774 177420 140780 177472
rect 140832 177460 140838 177472
rect 221550 177460 221556 177472
rect 140832 177432 221556 177460
rect 140832 177420 140838 177432
rect 221550 177420 221556 177432
rect 221608 177420 221614 177472
rect 238018 177420 238024 177472
rect 238076 177460 238082 177472
rect 353294 177460 353300 177472
rect 238076 177432 353300 177460
rect 238076 177420 238082 177432
rect 353294 177420 353300 177432
rect 353352 177420 353358 177472
rect 124214 177352 124220 177404
rect 124272 177392 124278 177404
rect 220078 177392 220084 177404
rect 124272 177364 220084 177392
rect 124272 177352 124278 177364
rect 220078 177352 220084 177364
rect 220136 177352 220142 177404
rect 240594 177352 240600 177404
rect 240652 177392 240658 177404
rect 394694 177392 394700 177404
rect 240652 177364 394700 177392
rect 240652 177352 240658 177364
rect 394694 177352 394700 177364
rect 394752 177352 394758 177404
rect 9674 177284 9680 177336
rect 9732 177324 9738 177336
rect 210326 177324 210332 177336
rect 9732 177296 210332 177324
rect 9732 177284 9738 177296
rect 210326 177284 210332 177296
rect 210384 177284 210390 177336
rect 211522 177284 211528 177336
rect 211580 177324 211586 177336
rect 226794 177324 226800 177336
rect 211580 177296 226800 177324
rect 211580 177284 211586 177296
rect 226794 177284 226800 177296
rect 226852 177284 226858 177336
rect 228266 177284 228272 177336
rect 228324 177324 228330 177336
rect 238018 177324 238024 177336
rect 228324 177296 238024 177324
rect 228324 177284 228330 177296
rect 238018 177284 238024 177296
rect 238076 177284 238082 177336
rect 249058 177284 249064 177336
rect 249116 177324 249122 177336
rect 496814 177324 496820 177336
rect 249116 177296 496820 177324
rect 249116 177284 249122 177296
rect 496814 177284 496820 177296
rect 496872 177284 496878 177336
rect 226886 176672 226892 176724
rect 226944 176712 226950 176724
rect 228174 176712 228180 176724
rect 226944 176684 228180 176712
rect 226944 176672 226950 176684
rect 228174 176672 228180 176684
rect 228232 176672 228238 176724
rect 31754 168988 31760 169040
rect 31812 169028 31818 169040
rect 203702 169028 203708 169040
rect 31812 169000 203708 169028
rect 31812 168988 31818 169000
rect 203702 168988 203708 169000
rect 203760 168988 203766 169040
rect 273990 166948 273996 167000
rect 274048 166988 274054 167000
rect 580166 166988 580172 167000
rect 274048 166960 580172 166988
rect 274048 166948 274054 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 196618 164200 196624 164212
rect 3384 164172 196624 164200
rect 3384 164160 3390 164172
rect 196618 164160 196624 164172
rect 196676 164160 196682 164212
rect 298922 153144 298928 153196
rect 298980 153184 298986 153196
rect 580166 153184 580172 153196
rect 298980 153156 580172 153184
rect 298980 153144 298986 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 192478 150396 192484 150408
rect 3384 150368 192484 150396
rect 3384 150356 3390 150368
rect 192478 150356 192484 150368
rect 192536 150356 192542 150408
rect 295978 139340 295984 139392
rect 296036 139380 296042 139392
rect 580166 139380 580172 139392
rect 296036 139352 580172 139380
rect 296036 139340 296042 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 268378 126896 268384 126948
rect 268436 126936 268442 126948
rect 580166 126936 580172 126948
rect 268436 126908 580172 126936
rect 268436 126896 268442 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 298830 113092 298836 113144
rect 298888 113132 298894 113144
rect 579798 113132 579804 113144
rect 298888 113104 579804 113132
rect 298888 113092 298894 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 199378 111772 199384 111784
rect 3200 111744 199384 111772
rect 3200 111732 3206 111744
rect 199378 111732 199384 111744
rect 199436 111732 199442 111784
rect 296070 100648 296076 100700
rect 296128 100688 296134 100700
rect 580166 100688 580172 100700
rect 296128 100660 580172 100688
rect 296128 100648 296134 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 232406 87796 232412 87848
rect 232464 87836 232470 87848
rect 288434 87836 288440 87848
rect 232464 87808 288440 87836
rect 232464 87796 232470 87808
rect 288434 87796 288440 87808
rect 288492 87796 288498 87848
rect 235258 87728 235264 87780
rect 235316 87768 235322 87780
rect 311894 87768 311900 87780
rect 235316 87740 311900 87768
rect 235316 87728 235322 87740
rect 311894 87728 311900 87740
rect 311952 87728 311958 87780
rect 239398 87660 239404 87712
rect 239456 87700 239462 87712
rect 375374 87700 375380 87712
rect 239456 87672 375380 87700
rect 239456 87660 239462 87672
rect 375374 87660 375380 87672
rect 375432 87660 375438 87712
rect 241882 87592 241888 87644
rect 241940 87632 241946 87644
rect 411254 87632 411260 87644
rect 241940 87604 411260 87632
rect 241940 87592 241946 87604
rect 411254 87592 411260 87604
rect 411312 87592 411318 87644
rect 265618 86912 265624 86964
rect 265676 86952 265682 86964
rect 580166 86952 580172 86964
rect 265676 86924 580172 86952
rect 265676 86912 265682 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 243538 86504 243544 86556
rect 243596 86544 243602 86556
rect 427814 86544 427820 86556
rect 243596 86516 427820 86544
rect 243596 86504 243602 86516
rect 427814 86504 427820 86516
rect 427872 86504 427878 86556
rect 244826 86436 244832 86488
rect 244884 86476 244890 86488
rect 447134 86476 447140 86488
rect 244884 86448 447140 86476
rect 244884 86436 244890 86448
rect 447134 86436 447140 86448
rect 447192 86436 447198 86488
rect 246206 86368 246212 86420
rect 246264 86408 246270 86420
rect 454034 86408 454040 86420
rect 246264 86380 454040 86408
rect 246264 86368 246270 86380
rect 454034 86368 454040 86380
rect 454092 86368 454098 86420
rect 247586 86300 247592 86352
rect 247644 86340 247650 86352
rect 478874 86340 478880 86352
rect 247644 86312 478880 86340
rect 247644 86300 247650 86312
rect 478874 86300 478880 86312
rect 478932 86300 478938 86352
rect 117314 86232 117320 86284
rect 117372 86272 117378 86284
rect 206278 86272 206284 86284
rect 117372 86244 206284 86272
rect 117372 86232 117378 86244
rect 206278 86232 206284 86244
rect 206336 86232 206342 86284
rect 250438 86232 250444 86284
rect 250496 86272 250502 86284
rect 517514 86272 517520 86284
rect 250496 86244 517520 86272
rect 250496 86232 250502 86244
rect 517514 86232 517520 86244
rect 517572 86232 517578 86284
rect 95234 83444 95240 83496
rect 95292 83484 95298 83496
rect 207842 83484 207848 83496
rect 95292 83456 207848 83484
rect 95292 83444 95298 83456
rect 207842 83444 207848 83456
rect 207900 83444 207906 83496
rect 244918 82220 244924 82272
rect 244976 82260 244982 82272
rect 365806 82260 365812 82272
rect 244976 82232 365812 82260
rect 244976 82220 244982 82232
rect 365806 82220 365812 82232
rect 365864 82220 365870 82272
rect 243446 82152 243452 82204
rect 243504 82192 243510 82204
rect 420914 82192 420920 82204
rect 243504 82164 420920 82192
rect 243504 82152 243510 82164
rect 420914 82152 420920 82164
rect 420972 82152 420978 82204
rect 278038 82084 278044 82136
rect 278096 82124 278102 82136
rect 581086 82124 581092 82136
rect 278096 82096 581092 82124
rect 278096 82084 278102 82096
rect 581086 82084 581092 82096
rect 581144 82084 581150 82136
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 200850 71720 200856 71732
rect 3476 71692 200856 71720
rect 3476 71680 3482 71692
rect 200850 71680 200856 71692
rect 200908 71680 200914 71732
rect 273898 60664 273904 60716
rect 273956 60704 273962 60716
rect 580166 60704 580172 60716
rect 273956 60676 580172 60704
rect 273956 60664 273962 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 256326 60052 256332 60104
rect 256384 60092 256390 60104
rect 400214 60092 400220 60104
rect 256384 60064 400220 60092
rect 256384 60052 256390 60064
rect 400214 60052 400220 60064
rect 400272 60052 400278 60104
rect 256234 59984 256240 60036
rect 256292 60024 256298 60036
rect 407114 60024 407120 60036
rect 256292 59996 407120 60024
rect 256292 59984 256298 59996
rect 407114 59984 407120 59996
rect 407172 59984 407178 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 79318 59344 79324 59356
rect 3108 59316 79324 59344
rect 3108 59304 3114 59316
rect 79318 59304 79324 59316
rect 79376 59304 79382 59356
rect 218606 46316 218612 46368
rect 218664 46356 218670 46368
rect 226610 46356 226616 46368
rect 218664 46328 226616 46356
rect 218664 46316 218670 46328
rect 226610 46316 226616 46328
rect 226668 46316 226674 46368
rect 162854 46248 162860 46300
rect 162912 46288 162918 46300
rect 222746 46288 222752 46300
rect 162912 46260 222752 46288
rect 162912 46248 162918 46260
rect 222746 46248 222752 46260
rect 222804 46248 222810 46300
rect 149054 46180 149060 46232
rect 149112 46220 149118 46232
rect 221458 46220 221464 46232
rect 149112 46192 221464 46220
rect 149112 46180 149118 46192
rect 221458 46180 221464 46192
rect 221516 46180 221522 46232
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 197998 33096 198004 33108
rect 3200 33068 198004 33096
rect 3200 33056 3206 33068
rect 197998 33056 198004 33068
rect 198056 33056 198062 33108
rect 298738 33056 298744 33108
rect 298796 33096 298802 33108
rect 580166 33096 580172 33108
rect 298796 33068 580172 33096
rect 298796 33056 298802 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 271138 31016 271144 31068
rect 271196 31056 271202 31068
rect 467834 31056 467840 31068
rect 271196 31028 467840 31056
rect 271196 31016 271202 31028
rect 467834 31016 467840 31028
rect 467892 31016 467898 31068
rect 269758 29588 269764 29640
rect 269816 29628 269822 29640
rect 460934 29628 460940 29640
rect 269816 29600 460940 29628
rect 269816 29588 269822 29600
rect 460934 29588 460940 29600
rect 460992 29588 460998 29640
rect 264238 28228 264244 28280
rect 264296 28268 264302 28280
rect 456886 28268 456892 28280
rect 264296 28240 456892 28268
rect 264296 28228 264302 28240
rect 456886 28228 456892 28240
rect 456944 28228 456950 28280
rect 237926 27208 237932 27260
rect 237984 27248 237990 27260
rect 350534 27248 350540 27260
rect 237984 27220 350540 27248
rect 237984 27208 237990 27220
rect 350534 27208 350540 27220
rect 350592 27208 350598 27260
rect 237834 27140 237840 27192
rect 237892 27180 237898 27192
rect 354674 27180 354680 27192
rect 237892 27152 354680 27180
rect 237892 27140 237898 27152
rect 354674 27140 354680 27152
rect 354732 27140 354738 27192
rect 239306 27072 239312 27124
rect 239364 27112 239370 27124
rect 368474 27112 368480 27124
rect 239364 27084 368480 27112
rect 239364 27072 239370 27084
rect 368474 27072 368480 27084
rect 368532 27072 368538 27124
rect 240502 27004 240508 27056
rect 240560 27044 240566 27056
rect 386414 27044 386420 27056
rect 240560 27016 386420 27044
rect 240560 27004 240566 27016
rect 386414 27004 386420 27016
rect 386472 27004 386478 27056
rect 240410 26936 240416 26988
rect 240468 26976 240474 26988
rect 397454 26976 397460 26988
rect 240468 26948 397460 26976
rect 240468 26936 240474 26948
rect 397454 26936 397460 26948
rect 397512 26936 397518 26988
rect 241790 26868 241796 26920
rect 241848 26908 241854 26920
rect 404354 26908 404360 26920
rect 241848 26880 404360 26908
rect 241848 26868 241854 26880
rect 404354 26868 404360 26880
rect 404412 26868 404418 26920
rect 232222 25916 232228 25968
rect 232280 25956 232286 25968
rect 280154 25956 280160 25968
rect 232280 25928 280160 25956
rect 232280 25916 232286 25928
rect 280154 25916 280160 25928
rect 280212 25916 280218 25968
rect 232314 25848 232320 25900
rect 232372 25888 232378 25900
rect 284386 25888 284392 25900
rect 232372 25860 284392 25888
rect 232372 25848 232378 25860
rect 284386 25848 284392 25860
rect 284444 25848 284450 25900
rect 232130 25780 232136 25832
rect 232188 25820 232194 25832
rect 287054 25820 287060 25832
rect 232188 25792 287060 25820
rect 232188 25780 232194 25792
rect 287054 25780 287060 25792
rect 287112 25780 287118 25832
rect 233786 25712 233792 25764
rect 233844 25752 233850 25764
rect 300854 25752 300860 25764
rect 233844 25724 300860 25752
rect 233844 25712 233850 25724
rect 300854 25712 300860 25724
rect 300912 25712 300918 25764
rect 235166 25644 235172 25696
rect 235224 25684 235230 25696
rect 318794 25684 318800 25696
rect 235224 25656 318800 25684
rect 235224 25644 235230 25656
rect 318794 25644 318800 25656
rect 318852 25644 318858 25696
rect 236454 25576 236460 25628
rect 236512 25616 236518 25628
rect 336734 25616 336740 25628
rect 236512 25588 336740 25616
rect 236512 25576 236518 25588
rect 336734 25576 336740 25588
rect 336792 25576 336798 25628
rect 255406 25508 255412 25560
rect 255464 25548 255470 25560
rect 578234 25548 578240 25560
rect 255464 25520 578240 25548
rect 255464 25508 255470 25520
rect 578234 25508 578240 25520
rect 578292 25508 578298 25560
rect 250346 24420 250352 24472
rect 250404 24460 250410 24472
rect 510614 24460 510620 24472
rect 250404 24432 510620 24460
rect 250404 24420 250410 24432
rect 510614 24420 510620 24432
rect 510672 24420 510678 24472
rect 250254 24352 250260 24404
rect 250312 24392 250318 24404
rect 514846 24392 514852 24404
rect 250312 24364 514852 24392
rect 250312 24352 250318 24364
rect 514846 24352 514852 24364
rect 514904 24352 514910 24404
rect 251726 24284 251732 24336
rect 251784 24324 251790 24336
rect 524414 24324 524420 24336
rect 251784 24296 524420 24324
rect 251784 24284 251790 24296
rect 524414 24284 524420 24296
rect 524472 24284 524478 24336
rect 251634 24216 251640 24268
rect 251692 24256 251698 24268
rect 528554 24256 528560 24268
rect 251692 24228 528560 24256
rect 251692 24216 251698 24228
rect 528554 24216 528560 24228
rect 528612 24216 528618 24268
rect 251542 24148 251548 24200
rect 251600 24188 251606 24200
rect 531314 24188 531320 24200
rect 251600 24160 531320 24188
rect 251600 24148 251606 24160
rect 531314 24148 531320 24160
rect 531372 24148 531378 24200
rect 254486 24080 254492 24132
rect 254544 24120 254550 24132
rect 567194 24120 567200 24132
rect 254544 24092 567200 24120
rect 254544 24080 254550 24092
rect 567194 24080 567200 24092
rect 567252 24080 567258 24132
rect 246022 23128 246028 23180
rect 246080 23168 246086 23180
rect 459554 23168 459560 23180
rect 246080 23140 459560 23168
rect 246080 23128 246086 23140
rect 459554 23128 459560 23140
rect 459612 23128 459618 23180
rect 246114 23060 246120 23112
rect 246172 23100 246178 23112
rect 463694 23100 463700 23112
rect 246172 23072 463700 23100
rect 246172 23060 246178 23072
rect 463694 23060 463700 23072
rect 463752 23060 463758 23112
rect 247494 22992 247500 23044
rect 247552 23032 247558 23044
rect 477494 23032 477500 23044
rect 247552 23004 477500 23032
rect 247552 22992 247558 23004
rect 477494 22992 477500 23004
rect 477552 22992 477558 23044
rect 247402 22924 247408 22976
rect 247460 22964 247466 22976
rect 481634 22964 481640 22976
rect 247460 22936 481640 22964
rect 247460 22924 247466 22936
rect 481634 22924 481640 22936
rect 481692 22924 481698 22976
rect 248874 22856 248880 22908
rect 248932 22896 248938 22908
rect 490006 22896 490012 22908
rect 248932 22868 490012 22896
rect 248932 22856 248938 22868
rect 490006 22856 490012 22868
rect 490064 22856 490070 22908
rect 248966 22788 248972 22840
rect 249024 22828 249030 22840
rect 492674 22828 492680 22840
rect 249024 22800 492680 22828
rect 249024 22788 249030 22800
rect 492674 22788 492680 22800
rect 492732 22788 492738 22840
rect 250162 22720 250168 22772
rect 250220 22760 250226 22772
rect 506566 22760 506572 22772
rect 250220 22732 506572 22760
rect 250220 22720 250226 22732
rect 506566 22720 506572 22732
rect 506624 22720 506630 22772
rect 240318 21632 240324 21684
rect 240376 21672 240382 21684
rect 396074 21672 396080 21684
rect 240376 21644 396080 21672
rect 240376 21632 240382 21644
rect 396074 21632 396080 21644
rect 396132 21632 396138 21684
rect 241698 21564 241704 21616
rect 241756 21604 241762 21616
rect 407206 21604 407212 21616
rect 241756 21576 407212 21604
rect 241756 21564 241762 21576
rect 407206 21564 407212 21576
rect 407264 21564 407270 21616
rect 244642 21496 244648 21548
rect 244700 21536 244706 21548
rect 438854 21536 438860 21548
rect 244700 21508 438860 21536
rect 244700 21496 244706 21508
rect 438854 21496 438860 21508
rect 438912 21496 438918 21548
rect 244458 21428 244464 21480
rect 244516 21468 244522 21480
rect 441614 21468 441620 21480
rect 244516 21440 441620 21468
rect 244516 21428 244522 21440
rect 441614 21428 441620 21440
rect 441672 21428 441678 21480
rect 244550 21360 244556 21412
rect 244608 21400 244614 21412
rect 448514 21400 448520 21412
rect 244608 21372 448520 21400
rect 244608 21360 244614 21372
rect 448514 21360 448520 21372
rect 448572 21360 448578 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 200758 20652 200764 20664
rect 3476 20624 200764 20652
rect 3476 20612 3482 20624
rect 200758 20612 200764 20624
rect 200816 20612 200822 20664
rect 235074 20272 235080 20324
rect 235132 20312 235138 20324
rect 317414 20312 317420 20324
rect 235132 20284 317420 20312
rect 235132 20272 235138 20284
rect 317414 20272 317420 20284
rect 317472 20272 317478 20324
rect 234982 20204 234988 20256
rect 235040 20244 235046 20256
rect 321554 20244 321560 20256
rect 235040 20216 321560 20244
rect 235040 20204 235046 20216
rect 321554 20204 321560 20216
rect 321612 20204 321618 20256
rect 237742 20136 237748 20188
rect 237800 20176 237806 20188
rect 349154 20176 349160 20188
rect 237800 20148 349160 20176
rect 237800 20136 237806 20148
rect 349154 20136 349160 20148
rect 349212 20136 349218 20188
rect 239122 20068 239128 20120
rect 239180 20108 239186 20120
rect 367094 20108 367100 20120
rect 239180 20080 367100 20108
rect 239180 20068 239186 20080
rect 367094 20068 367100 20080
rect 367152 20068 367158 20120
rect 239030 20000 239036 20052
rect 239088 20040 239094 20052
rect 371234 20040 371240 20052
rect 239088 20012 371240 20040
rect 239088 20000 239094 20012
rect 371234 20000 371240 20012
rect 371292 20000 371298 20052
rect 239214 19932 239220 19984
rect 239272 19972 239278 19984
rect 373994 19972 374000 19984
rect 239272 19944 374000 19972
rect 239272 19932 239278 19944
rect 373994 19932 374000 19944
rect 374052 19932 374058 19984
rect 232038 18912 232044 18964
rect 232096 18952 232102 18964
rect 285674 18952 285680 18964
rect 232096 18924 285680 18952
rect 232096 18912 232102 18924
rect 285674 18912 285680 18924
rect 285732 18912 285738 18964
rect 233602 18844 233608 18896
rect 233660 18884 233666 18896
rect 296714 18884 296720 18896
rect 233660 18856 296720 18884
rect 233660 18844 233666 18856
rect 296714 18844 296720 18856
rect 296772 18844 296778 18896
rect 233694 18776 233700 18828
rect 233752 18816 233758 18828
rect 299566 18816 299572 18828
rect 233752 18788 299572 18816
rect 233752 18776 233758 18788
rect 299566 18776 299572 18788
rect 299624 18776 299630 18828
rect 233510 18708 233516 18760
rect 233568 18748 233574 18760
rect 303614 18748 303620 18760
rect 233568 18720 303620 18748
rect 233568 18708 233574 18720
rect 303614 18708 303620 18720
rect 303672 18708 303678 18760
rect 234890 18640 234896 18692
rect 234948 18680 234954 18692
rect 314654 18680 314660 18692
rect 234948 18652 314660 18680
rect 234948 18640 234954 18652
rect 314654 18640 314660 18652
rect 314712 18640 314718 18692
rect 247310 18572 247316 18624
rect 247368 18612 247374 18624
rect 471974 18612 471980 18624
rect 247368 18584 471980 18612
rect 247368 18572 247374 18584
rect 471974 18572 471980 18584
rect 472032 18572 472038 18624
rect 233878 17620 233884 17672
rect 233936 17660 233942 17672
rect 271874 17660 271880 17672
rect 233936 17632 271880 17660
rect 233936 17620 233942 17632
rect 271874 17620 271880 17632
rect 271932 17620 271938 17672
rect 231946 17552 231952 17604
rect 232004 17592 232010 17604
rect 278774 17592 278780 17604
rect 232004 17564 278780 17592
rect 232004 17552 232010 17564
rect 278774 17552 278780 17564
rect 278832 17552 278838 17604
rect 231854 17484 231860 17536
rect 231912 17524 231918 17536
rect 282914 17524 282920 17536
rect 231912 17496 282920 17524
rect 231912 17484 231918 17496
rect 282914 17484 282920 17496
rect 282972 17484 282978 17536
rect 240226 17416 240232 17468
rect 240284 17456 240290 17468
rect 389174 17456 389180 17468
rect 240284 17428 389180 17456
rect 240284 17416 240290 17428
rect 389174 17416 389180 17428
rect 389232 17416 389238 17468
rect 254394 17348 254400 17400
rect 254452 17388 254458 17400
rect 563054 17388 563060 17400
rect 254452 17360 563060 17388
rect 254452 17348 254458 17360
rect 563054 17348 563060 17360
rect 563112 17348 563118 17400
rect 254210 17280 254216 17332
rect 254268 17320 254274 17332
rect 565814 17320 565820 17332
rect 254268 17292 565820 17320
rect 254268 17280 254274 17292
rect 565814 17280 565820 17292
rect 565872 17280 565878 17332
rect 254302 17212 254308 17264
rect 254360 17252 254366 17264
rect 569954 17252 569960 17264
rect 254360 17224 569960 17252
rect 254360 17212 254366 17224
rect 569954 17212 569960 17224
rect 570012 17212 570018 17264
rect 251450 16124 251456 16176
rect 251508 16164 251514 16176
rect 527818 16164 527824 16176
rect 251508 16136 527824 16164
rect 251508 16124 251514 16136
rect 527818 16124 527824 16136
rect 527876 16124 527882 16176
rect 251358 16056 251364 16108
rect 251416 16096 251422 16108
rect 531406 16096 531412 16108
rect 251416 16068 531412 16096
rect 251416 16056 251422 16068
rect 531406 16056 531412 16068
rect 531464 16056 531470 16108
rect 253106 15988 253112 16040
rect 253164 16028 253170 16040
rect 545482 16028 545488 16040
rect 253164 16000 545488 16028
rect 253164 15988 253170 16000
rect 545482 15988 545488 16000
rect 545540 15988 545546 16040
rect 114002 15920 114008 15972
rect 114060 15960 114066 15972
rect 218514 15960 218520 15972
rect 114060 15932 218520 15960
rect 114060 15920 114066 15932
rect 218514 15920 218520 15932
rect 218572 15920 218578 15972
rect 253014 15920 253020 15972
rect 253072 15960 253078 15972
rect 548610 15960 548616 15972
rect 253072 15932 548616 15960
rect 253072 15920 253078 15932
rect 548610 15920 548616 15932
rect 548668 15920 548674 15972
rect 35986 15852 35992 15904
rect 36044 15892 36050 15904
rect 212902 15892 212908 15904
rect 36044 15864 212908 15892
rect 36044 15852 36050 15864
rect 212902 15852 212908 15864
rect 212960 15852 212966 15904
rect 252922 15852 252928 15904
rect 252980 15892 252986 15904
rect 552658 15892 552664 15904
rect 252980 15864 552664 15892
rect 252980 15852 252986 15864
rect 552658 15852 552664 15864
rect 552716 15852 552722 15904
rect 123018 14900 123024 14952
rect 123076 14940 123082 14952
rect 219986 14940 219992 14952
rect 123076 14912 219992 14940
rect 123076 14900 123082 14912
rect 219986 14900 219992 14912
rect 220044 14900 220050 14952
rect 256142 14900 256148 14952
rect 256200 14940 256206 14952
rect 422570 14940 422576 14952
rect 256200 14912 422576 14940
rect 256200 14900 256206 14912
rect 422570 14900 422576 14912
rect 422628 14900 422634 14952
rect 105722 14832 105728 14884
rect 105780 14872 105786 14884
rect 218422 14872 218428 14884
rect 105780 14844 218428 14872
rect 105780 14832 105786 14844
rect 218422 14832 218428 14844
rect 218480 14832 218486 14884
rect 248598 14832 248604 14884
rect 248656 14872 248662 14884
rect 492306 14872 492312 14884
rect 248656 14844 492312 14872
rect 248656 14832 248662 14844
rect 492306 14832 492312 14844
rect 492364 14832 492370 14884
rect 98178 14764 98184 14816
rect 98236 14804 98242 14816
rect 216950 14804 216956 14816
rect 98236 14776 216956 14804
rect 98236 14764 98242 14776
rect 216950 14764 216956 14776
rect 217008 14764 217014 14816
rect 248782 14764 248788 14816
rect 248840 14804 248846 14816
rect 495434 14804 495440 14816
rect 248840 14776 495440 14804
rect 248840 14764 248846 14776
rect 495434 14764 495440 14776
rect 495492 14764 495498 14816
rect 74994 14696 75000 14748
rect 75052 14736 75058 14748
rect 215938 14736 215944 14748
rect 75052 14708 215944 14736
rect 75052 14696 75058 14708
rect 215938 14696 215944 14708
rect 215996 14696 216002 14748
rect 248506 14696 248512 14748
rect 248564 14736 248570 14748
rect 498930 14736 498936 14748
rect 248564 14708 498936 14736
rect 248564 14696 248570 14708
rect 498930 14696 498936 14708
rect 498988 14696 498994 14748
rect 44174 14628 44180 14680
rect 44232 14668 44238 14680
rect 212810 14668 212816 14680
rect 44232 14640 212816 14668
rect 44232 14628 44238 14640
rect 212810 14628 212816 14640
rect 212868 14628 212874 14680
rect 248690 14628 248696 14680
rect 248748 14668 248754 14680
rect 502978 14668 502984 14680
rect 248748 14640 502984 14668
rect 248748 14628 248754 14640
rect 502978 14628 502984 14640
rect 503036 14628 503042 14680
rect 34514 14560 34520 14612
rect 34572 14600 34578 14612
rect 211798 14600 211804 14612
rect 34572 14572 211804 14600
rect 34572 14560 34578 14572
rect 211798 14560 211804 14572
rect 211856 14560 211862 14612
rect 250070 14560 250076 14612
rect 250128 14600 250134 14612
rect 509602 14600 509608 14612
rect 250128 14572 509608 14600
rect 250128 14560 250134 14572
rect 509602 14560 509608 14572
rect 509660 14560 509666 14612
rect 22554 14492 22560 14544
rect 22612 14532 22618 14544
rect 211430 14532 211436 14544
rect 22612 14504 211436 14532
rect 22612 14492 22618 14504
rect 211430 14492 211436 14504
rect 211488 14492 211494 14544
rect 249978 14492 249984 14544
rect 250036 14532 250042 14544
rect 513374 14532 513380 14544
rect 250036 14504 513380 14532
rect 250036 14492 250042 14504
rect 513374 14492 513380 14504
rect 513432 14492 513438 14544
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 211338 14464 211344 14476
rect 18012 14436 211344 14464
rect 18012 14424 18018 14436
rect 211338 14424 211344 14436
rect 211396 14424 211402 14476
rect 249886 14424 249892 14476
rect 249944 14464 249950 14476
rect 517146 14464 517152 14476
rect 249944 14436 517152 14464
rect 249944 14424 249950 14436
rect 517146 14424 517152 14436
rect 517204 14424 517210 14476
rect 80882 13540 80888 13592
rect 80940 13580 80946 13592
rect 215846 13580 215852 13592
rect 80940 13552 215852 13580
rect 80940 13540 80946 13552
rect 215846 13540 215852 13552
rect 215904 13540 215910 13592
rect 77386 13472 77392 13524
rect 77444 13512 77450 13524
rect 215570 13512 215576 13524
rect 77444 13484 215576 13512
rect 77444 13472 77450 13484
rect 215570 13472 215576 13484
rect 215628 13472 215634 13524
rect 243354 13472 243360 13524
rect 243412 13512 243418 13524
rect 425698 13512 425704 13524
rect 243412 13484 425704 13512
rect 243412 13472 243418 13484
rect 425698 13472 425704 13484
rect 425756 13472 425762 13524
rect 73338 13404 73344 13456
rect 73396 13444 73402 13456
rect 215662 13444 215668 13456
rect 73396 13416 215668 13444
rect 73396 13404 73402 13416
rect 215662 13404 215668 13416
rect 215720 13404 215726 13456
rect 245930 13404 245936 13456
rect 245988 13444 245994 13456
rect 459186 13444 459192 13456
rect 245988 13416 459192 13444
rect 245988 13404 245994 13416
rect 459186 13404 459192 13416
rect 459244 13404 459250 13456
rect 69842 13336 69848 13388
rect 69900 13376 69906 13388
rect 215754 13376 215760 13388
rect 69900 13348 215760 13376
rect 69900 13336 69906 13348
rect 215754 13336 215760 13348
rect 215812 13336 215818 13388
rect 245746 13336 245752 13388
rect 245804 13376 245810 13388
rect 462314 13376 462320 13388
rect 245804 13348 462320 13376
rect 245804 13336 245810 13348
rect 462314 13336 462320 13348
rect 462372 13336 462378 13388
rect 59354 13268 59360 13320
rect 59412 13308 59418 13320
rect 214374 13308 214380 13320
rect 59412 13280 214380 13308
rect 59412 13268 59418 13280
rect 214374 13268 214380 13280
rect 214432 13268 214438 13320
rect 245838 13268 245844 13320
rect 245896 13308 245902 13320
rect 465810 13308 465816 13320
rect 245896 13280 465816 13308
rect 245896 13268 245902 13280
rect 465810 13268 465816 13280
rect 465868 13268 465874 13320
rect 56042 13200 56048 13252
rect 56100 13240 56106 13252
rect 214282 13240 214288 13252
rect 56100 13212 214288 13240
rect 56100 13200 56106 13212
rect 214282 13200 214288 13212
rect 214340 13200 214346 13252
rect 247034 13200 247040 13252
rect 247092 13240 247098 13252
rect 473446 13240 473452 13252
rect 247092 13212 473452 13240
rect 247092 13200 247098 13212
rect 473446 13200 473452 13212
rect 473504 13200 473510 13252
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 210234 13172 210240 13184
rect 8812 13144 210240 13172
rect 8812 13132 8818 13144
rect 210234 13132 210240 13144
rect 210292 13132 210298 13184
rect 247218 13132 247224 13184
rect 247276 13172 247282 13184
rect 476482 13172 476488 13184
rect 247276 13144 476488 13172
rect 247276 13132 247282 13144
rect 476482 13132 476488 13144
rect 476540 13132 476546 13184
rect 3602 13064 3608 13116
rect 3660 13104 3666 13116
rect 210142 13104 210148 13116
rect 3660 13076 210148 13104
rect 3660 13064 3666 13076
rect 210142 13064 210148 13076
rect 210200 13064 210206 13116
rect 247126 13064 247132 13116
rect 247184 13104 247190 13116
rect 481726 13104 481732 13116
rect 247184 13076 481732 13104
rect 247184 13064 247190 13076
rect 481726 13064 481732 13076
rect 481784 13064 481790 13116
rect 240134 12112 240140 12164
rect 240192 12152 240198 12164
rect 390646 12152 390652 12164
rect 240192 12124 390652 12152
rect 240192 12112 240198 12124
rect 390646 12112 390652 12124
rect 390704 12112 390710 12164
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 178678 12084 178684 12096
rect 15988 12056 178684 12084
rect 15988 12044 15994 12056
rect 178678 12044 178684 12056
rect 178736 12044 178742 12096
rect 178770 12044 178776 12096
rect 178828 12084 178834 12096
rect 214190 12084 214196 12096
rect 178828 12056 214196 12084
rect 178828 12044 178834 12056
rect 214190 12044 214196 12056
rect 214248 12044 214254 12096
rect 243262 12044 243268 12096
rect 243320 12084 243326 12096
rect 423766 12084 423772 12096
rect 243320 12056 423772 12084
rect 243320 12044 243326 12056
rect 423766 12044 423772 12056
rect 423824 12044 423830 12096
rect 44266 11976 44272 12028
rect 44324 12016 44330 12028
rect 213270 12016 213276 12028
rect 44324 11988 213276 12016
rect 44324 11976 44330 11988
rect 213270 11976 213276 11988
rect 213328 11976 213334 12028
rect 243078 11976 243084 12028
rect 243136 12016 243142 12028
rect 426802 12016 426808 12028
rect 243136 11988 426808 12016
rect 243136 11976 243142 11988
rect 426802 11976 426808 11988
rect 426860 11976 426866 12028
rect 36722 11908 36728 11960
rect 36780 11948 36786 11960
rect 212626 11948 212632 11960
rect 36780 11920 212632 11948
rect 36780 11908 36786 11920
rect 212626 11908 212632 11920
rect 212684 11908 212690 11960
rect 243170 11908 243176 11960
rect 243228 11948 243234 11960
rect 430850 11948 430856 11960
rect 243228 11920 430856 11948
rect 243228 11908 243234 11920
rect 430850 11908 430856 11920
rect 430908 11908 430914 11960
rect 33594 11840 33600 11892
rect 33652 11880 33658 11892
rect 212718 11880 212724 11892
rect 33652 11852 212724 11880
rect 33652 11840 33658 11852
rect 212718 11840 212724 11852
rect 212776 11840 212782 11892
rect 244274 11840 244280 11892
rect 244332 11880 244338 11892
rect 445018 11880 445024 11892
rect 244332 11852 445024 11880
rect 244332 11840 244338 11852
rect 445018 11840 445024 11852
rect 445076 11840 445082 11892
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 211614 11812 211620 11824
rect 26292 11784 211620 11812
rect 26292 11772 26298 11784
rect 211614 11772 211620 11784
rect 211672 11772 211678 11824
rect 244366 11772 244372 11824
rect 244424 11812 244430 11824
rect 448606 11812 448612 11824
rect 244424 11784 448612 11812
rect 244424 11772 244430 11784
rect 448606 11772 448612 11784
rect 448664 11772 448670 11824
rect 21818 11704 21824 11756
rect 21876 11744 21882 11756
rect 212350 11744 212356 11756
rect 21876 11716 212356 11744
rect 21876 11704 21882 11716
rect 212350 11704 212356 11716
rect 212408 11704 212414 11756
rect 245654 11704 245660 11756
rect 245712 11744 245718 11756
rect 455690 11744 455696 11756
rect 245712 11716 455696 11744
rect 245712 11704 245718 11716
rect 455690 11704 455696 11716
rect 455748 11704 455754 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 171778 10752 171784 10804
rect 171836 10792 171842 10804
rect 218330 10792 218336 10804
rect 171836 10764 218336 10792
rect 171836 10752 171842 10764
rect 218330 10752 218336 10764
rect 218388 10752 218394 10804
rect 111610 10684 111616 10736
rect 111668 10724 111674 10736
rect 218698 10724 218704 10736
rect 111668 10696 218704 10724
rect 111668 10684 111674 10696
rect 218698 10684 218704 10696
rect 218756 10684 218762 10736
rect 108114 10616 108120 10668
rect 108172 10656 108178 10668
rect 218790 10656 218796 10668
rect 108172 10628 218796 10656
rect 108172 10616 108178 10628
rect 218790 10616 218796 10628
rect 218848 10616 218854 10668
rect 238846 10616 238852 10668
rect 238904 10656 238910 10668
rect 374086 10656 374092 10668
rect 238904 10628 374092 10656
rect 238904 10616 238910 10628
rect 374086 10616 374092 10628
rect 374144 10616 374150 10668
rect 104066 10548 104072 10600
rect 104124 10588 104130 10600
rect 218238 10588 218244 10600
rect 104124 10560 218244 10588
rect 104124 10548 104130 10560
rect 218238 10548 218244 10560
rect 218296 10548 218302 10600
rect 247678 10548 247684 10600
rect 247736 10588 247742 10600
rect 384298 10588 384304 10600
rect 247736 10560 384304 10588
rect 247736 10548 247742 10560
rect 384298 10548 384304 10560
rect 384356 10548 384362 10600
rect 97442 10480 97448 10532
rect 97500 10520 97506 10532
rect 216766 10520 216772 10532
rect 97500 10492 216772 10520
rect 97500 10480 97506 10492
rect 216766 10480 216772 10492
rect 216824 10480 216830 10532
rect 242434 10480 242440 10532
rect 242492 10520 242498 10532
rect 379514 10520 379520 10532
rect 242492 10492 379520 10520
rect 242492 10480 242498 10492
rect 379514 10480 379520 10492
rect 379572 10480 379578 10532
rect 93946 10412 93952 10464
rect 94004 10452 94010 10464
rect 216858 10452 216864 10464
rect 94004 10424 216864 10452
rect 94004 10412 94010 10424
rect 216858 10412 216864 10424
rect 216916 10412 216922 10464
rect 238938 10412 238944 10464
rect 238996 10452 239002 10464
rect 377674 10452 377680 10464
rect 238996 10424 377680 10452
rect 238996 10412 239002 10424
rect 377674 10412 377680 10424
rect 377732 10412 377738 10464
rect 89898 10344 89904 10396
rect 89956 10384 89962 10396
rect 217410 10384 217416 10396
rect 89956 10356 217416 10384
rect 89956 10344 89962 10356
rect 217410 10344 217416 10356
rect 217468 10344 217474 10396
rect 241514 10344 241520 10396
rect 241572 10384 241578 10396
rect 406010 10384 406016 10396
rect 241572 10356 406016 10384
rect 241572 10344 241578 10356
rect 406010 10344 406016 10356
rect 406068 10344 406074 10396
rect 11146 10276 11152 10328
rect 11204 10316 11210 10328
rect 188338 10316 188344 10328
rect 11204 10288 188344 10316
rect 11204 10276 11210 10288
rect 188338 10276 188344 10288
rect 188396 10276 188402 10328
rect 241606 10276 241612 10328
rect 241664 10316 241670 10328
rect 409138 10316 409144 10328
rect 241664 10288 409144 10316
rect 241664 10276 241670 10288
rect 409138 10276 409144 10288
rect 409196 10276 409202 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 79686 9324 79692 9376
rect 79744 9364 79750 9376
rect 216122 9364 216128 9376
rect 79744 9336 216128 9364
rect 79744 9324 79750 9336
rect 216122 9324 216128 9336
rect 216180 9324 216186 9376
rect 76190 9256 76196 9308
rect 76248 9296 76254 9308
rect 215478 9296 215484 9308
rect 76248 9268 215484 9296
rect 76248 9256 76254 9268
rect 215478 9256 215484 9268
rect 215536 9256 215542 9308
rect 237650 9256 237656 9308
rect 237708 9296 237714 9308
rect 349246 9296 349252 9308
rect 237708 9268 349252 9296
rect 237708 9256 237714 9268
rect 349246 9256 349252 9268
rect 349304 9256 349310 9308
rect 72602 9188 72608 9240
rect 72660 9228 72666 9240
rect 216214 9228 216220 9240
rect 72660 9200 216220 9228
rect 72660 9188 72666 9200
rect 216214 9188 216220 9200
rect 216272 9188 216278 9240
rect 237558 9188 237564 9240
rect 237616 9228 237622 9240
rect 352834 9228 352840 9240
rect 237616 9200 352840 9228
rect 237616 9188 237622 9200
rect 352834 9188 352840 9200
rect 352892 9188 352898 9240
rect 62022 9120 62028 9172
rect 62080 9160 62086 9172
rect 214098 9160 214104 9172
rect 62080 9132 214104 9160
rect 62080 9120 62086 9132
rect 214098 9120 214104 9132
rect 214156 9120 214162 9172
rect 237466 9120 237472 9172
rect 237524 9160 237530 9172
rect 356330 9160 356336 9172
rect 237524 9132 356336 9160
rect 237524 9120 237530 9132
rect 356330 9120 356336 9132
rect 356388 9120 356394 9172
rect 58434 9052 58440 9104
rect 58492 9092 58498 9104
rect 214006 9092 214012 9104
rect 58492 9064 214012 9092
rect 58492 9052 58498 9064
rect 214006 9052 214012 9064
rect 214064 9052 214070 9104
rect 237374 9052 237380 9104
rect 237432 9092 237438 9104
rect 359918 9092 359924 9104
rect 237432 9064 359924 9092
rect 237432 9052 237438 9064
rect 359918 9052 359924 9064
rect 359976 9052 359982 9104
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 210050 9024 210056 9036
rect 7708 8996 210056 9024
rect 7708 8984 7714 8996
rect 210050 8984 210056 8996
rect 210108 8984 210114 9036
rect 238754 8984 238760 9036
rect 238812 9024 238818 9036
rect 370590 9024 370596 9036
rect 238812 8996 370596 9024
rect 238812 8984 238818 8996
rect 370590 8984 370596 8996
rect 370648 8984 370654 9036
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 209958 8956 209964 8968
rect 2924 8928 209964 8956
rect 2924 8916 2930 8928
rect 209958 8916 209964 8928
rect 210016 8916 210022 8968
rect 257430 8916 257436 8968
rect 257488 8956 257494 8968
rect 415486 8956 415492 8968
rect 257488 8928 415492 8956
rect 257488 8916 257494 8928
rect 415486 8916 415492 8928
rect 415544 8916 415550 8968
rect 197906 7964 197912 8016
rect 197964 8004 197970 8016
rect 225414 8004 225420 8016
rect 197964 7976 225420 8004
rect 197964 7964 197970 7976
rect 225414 7964 225420 7976
rect 225472 7964 225478 8016
rect 158898 7896 158904 7948
rect 158956 7936 158962 7948
rect 222654 7936 222660 7948
rect 158956 7908 222660 7936
rect 158956 7896 158962 7908
rect 222654 7896 222660 7908
rect 222712 7896 222718 7948
rect 151906 7828 151912 7880
rect 151964 7868 151970 7880
rect 221090 7868 221096 7880
rect 151964 7840 221096 7868
rect 151964 7828 151970 7840
rect 221090 7828 221096 7840
rect 221148 7828 221154 7880
rect 148318 7760 148324 7812
rect 148376 7800 148382 7812
rect 221182 7800 221188 7812
rect 148376 7772 221188 7800
rect 148376 7760 148382 7772
rect 221182 7760 221188 7772
rect 221240 7760 221246 7812
rect 233418 7760 233424 7812
rect 233476 7800 233482 7812
rect 306742 7800 306748 7812
rect 233476 7772 306748 7800
rect 233476 7760 233482 7772
rect 306742 7760 306748 7772
rect 306800 7760 306806 7812
rect 144730 7692 144736 7744
rect 144788 7732 144794 7744
rect 221274 7732 221280 7744
rect 144788 7704 221280 7732
rect 144788 7692 144794 7704
rect 221274 7692 221280 7704
rect 221332 7692 221338 7744
rect 234706 7692 234712 7744
rect 234764 7732 234770 7744
rect 320910 7732 320916 7744
rect 234764 7704 320916 7732
rect 234764 7692 234770 7704
rect 320910 7692 320916 7704
rect 320968 7692 320974 7744
rect 142430 7624 142436 7676
rect 142488 7664 142494 7676
rect 221366 7664 221372 7676
rect 142488 7636 221372 7664
rect 142488 7624 142494 7636
rect 221366 7624 221372 7636
rect 221424 7624 221430 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 324406 7664 324412 7676
rect 234856 7636 324412 7664
rect 234856 7624 234862 7636
rect 324406 7624 324412 7636
rect 324464 7624 324470 7676
rect 54938 7556 54944 7608
rect 54996 7596 55002 7608
rect 214742 7596 214748 7608
rect 54996 7568 214748 7596
rect 54996 7556 55002 7568
rect 214742 7556 214748 7568
rect 214800 7556 214806 7608
rect 252830 7556 252836 7608
rect 252888 7596 252894 7608
rect 553762 7596 553768 7608
rect 252888 7568 553768 7596
rect 252888 7556 252894 7568
rect 553762 7556 553768 7568
rect 553820 7556 553826 7608
rect 230750 6808 230756 6860
rect 230808 6848 230814 6860
rect 267734 6848 267740 6860
rect 230808 6820 267740 6848
rect 230808 6808 230814 6820
rect 267734 6808 267740 6820
rect 267792 6808 267798 6860
rect 230658 6740 230664 6792
rect 230716 6780 230722 6792
rect 268838 6780 268844 6792
rect 230716 6752 268844 6780
rect 230716 6740 230722 6752
rect 268838 6740 268844 6752
rect 268896 6740 268902 6792
rect 234614 6672 234620 6724
rect 234672 6712 234678 6724
rect 317322 6712 317328 6724
rect 234672 6684 317328 6712
rect 234672 6672 234678 6684
rect 317322 6672 317328 6684
rect 317380 6672 317386 6724
rect 200298 6604 200304 6656
rect 200356 6644 200362 6656
rect 225322 6644 225328 6656
rect 200356 6616 225328 6644
rect 200356 6604 200362 6616
rect 225322 6604 225328 6616
rect 225380 6604 225386 6656
rect 236270 6604 236276 6656
rect 236328 6644 236334 6656
rect 332686 6644 332692 6656
rect 236328 6616 332692 6644
rect 236328 6604 236334 6616
rect 332686 6604 332692 6616
rect 332744 6604 332750 6656
rect 187326 6536 187332 6588
rect 187384 6576 187390 6588
rect 223850 6576 223856 6588
rect 187384 6548 223856 6576
rect 187384 6536 187390 6548
rect 223850 6536 223856 6548
rect 223908 6536 223914 6588
rect 236178 6536 236184 6588
rect 236236 6576 236242 6588
rect 336274 6576 336280 6588
rect 236236 6548 336280 6576
rect 236236 6536 236242 6548
rect 336274 6536 336280 6548
rect 336332 6536 336338 6588
rect 183738 6468 183744 6520
rect 183796 6508 183802 6520
rect 223758 6508 223764 6520
rect 183796 6480 223764 6508
rect 183796 6468 183802 6480
rect 223758 6468 223764 6480
rect 223816 6468 223822 6520
rect 236362 6468 236368 6520
rect 236420 6508 236426 6520
rect 342162 6508 342168 6520
rect 236420 6480 342168 6508
rect 236420 6468 236426 6480
rect 342162 6468 342168 6480
rect 342220 6468 342226 6520
rect 180242 6400 180248 6452
rect 180300 6440 180306 6452
rect 224034 6440 224040 6452
rect 180300 6412 224040 6440
rect 180300 6400 180306 6412
rect 224034 6400 224040 6412
rect 224092 6400 224098 6452
rect 242894 6400 242900 6452
rect 242952 6440 242958 6452
rect 418982 6440 418988 6452
rect 242952 6412 418988 6440
rect 242952 6400 242958 6412
rect 418982 6400 418988 6412
rect 419040 6400 419046 6452
rect 176746 6332 176752 6384
rect 176804 6372 176810 6384
rect 223942 6372 223948 6384
rect 176804 6344 223948 6372
rect 176804 6332 176810 6344
rect 223942 6332 223948 6344
rect 224000 6332 224006 6384
rect 242986 6332 242992 6384
rect 243044 6372 243050 6384
rect 420178 6372 420184 6384
rect 243044 6344 420184 6372
rect 243044 6332 243050 6344
rect 420178 6332 420184 6344
rect 420236 6332 420242 6384
rect 169570 6264 169576 6316
rect 169628 6304 169634 6316
rect 222562 6304 222568 6316
rect 169628 6276 222568 6304
rect 169628 6264 169634 6276
rect 222562 6264 222568 6276
rect 222620 6264 222626 6316
rect 256050 6264 256056 6316
rect 256108 6304 256114 6316
rect 562042 6304 562048 6316
rect 256108 6276 562048 6304
rect 256108 6264 256114 6276
rect 562042 6264 562048 6276
rect 562100 6264 562106 6316
rect 134150 6196 134156 6248
rect 134208 6236 134214 6248
rect 219894 6236 219900 6248
rect 134208 6208 219900 6236
rect 134208 6196 134214 6208
rect 219894 6196 219900 6208
rect 219952 6196 219958 6248
rect 254118 6196 254124 6248
rect 254176 6236 254182 6248
rect 569126 6236 569132 6248
rect 254176 6208 569132 6236
rect 254176 6196 254182 6208
rect 569126 6196 569132 6208
rect 569184 6196 569190 6248
rect 128170 6128 128176 6180
rect 128228 6168 128234 6180
rect 219802 6168 219808 6180
rect 128228 6140 219808 6168
rect 128228 6128 128234 6140
rect 219802 6128 219808 6140
rect 219860 6128 219866 6180
rect 254026 6128 254032 6180
rect 254084 6168 254090 6180
rect 572714 6168 572720 6180
rect 254084 6140 572720 6168
rect 254084 6128 254090 6140
rect 572714 6128 572720 6140
rect 572772 6128 572778 6180
rect 230934 6060 230940 6112
rect 230992 6100 230998 6112
rect 265342 6100 265348 6112
rect 230992 6072 265348 6100
rect 230992 6060 230998 6072
rect 265342 6060 265348 6072
rect 265400 6060 265406 6112
rect 230842 5992 230848 6044
rect 230900 6032 230906 6044
rect 261754 6032 261760 6044
rect 230900 6004 261760 6032
rect 230900 5992 230906 6004
rect 261754 5992 261760 6004
rect 261812 5992 261818 6044
rect 201586 5380 201592 5432
rect 201644 5420 201650 5432
rect 225782 5420 225788 5432
rect 201644 5392 225788 5420
rect 201644 5380 201650 5392
rect 225782 5380 225788 5392
rect 225840 5380 225846 5432
rect 196802 5312 196808 5364
rect 196860 5352 196866 5364
rect 225874 5352 225880 5364
rect 196860 5324 225880 5352
rect 196860 5312 196866 5324
rect 225874 5312 225880 5324
rect 225932 5312 225938 5364
rect 166074 5244 166080 5296
rect 166132 5284 166138 5296
rect 222378 5284 222384 5296
rect 166132 5256 222384 5284
rect 166132 5244 166138 5256
rect 222378 5244 222384 5256
rect 222436 5244 222442 5296
rect 150618 5176 150624 5228
rect 150676 5216 150682 5228
rect 150676 5188 156736 5216
rect 150676 5176 150682 5188
rect 147122 5108 147128 5160
rect 147180 5148 147186 5160
rect 147180 5120 156552 5148
rect 147180 5108 147186 5120
rect 156524 5012 156552 5120
rect 156708 5080 156736 5188
rect 162486 5176 162492 5228
rect 162544 5216 162550 5228
rect 222470 5216 222476 5228
rect 162544 5188 222476 5216
rect 162544 5176 162550 5188
rect 222470 5176 222476 5188
rect 222528 5176 222534 5228
rect 249794 5176 249800 5228
rect 249852 5216 249858 5228
rect 519538 5216 519544 5228
rect 249852 5188 519544 5216
rect 249852 5176 249858 5188
rect 519538 5176 519544 5188
rect 519596 5176 519602 5228
rect 157794 5108 157800 5160
rect 157852 5148 157858 5160
rect 223206 5148 223212 5160
rect 157852 5120 223212 5148
rect 157852 5108 157858 5120
rect 223206 5108 223212 5120
rect 223264 5108 223270 5160
rect 251174 5108 251180 5160
rect 251232 5148 251238 5160
rect 533706 5148 533712 5160
rect 251232 5120 533712 5148
rect 251232 5108 251238 5120
rect 533706 5108 533712 5120
rect 533764 5108 533770 5160
rect 221642 5080 221648 5092
rect 156708 5052 221648 5080
rect 221642 5040 221648 5052
rect 221700 5040 221706 5092
rect 251266 5040 251272 5092
rect 251324 5080 251330 5092
rect 537202 5080 537208 5092
rect 251324 5052 537208 5080
rect 251324 5040 251330 5052
rect 537202 5040 537208 5052
rect 537260 5040 537266 5092
rect 220906 5012 220912 5024
rect 156524 4984 220912 5012
rect 220906 4972 220912 4984
rect 220964 4972 220970 5024
rect 252646 4972 252652 5024
rect 252704 5012 252710 5024
rect 547874 5012 547880 5024
rect 252704 4984 547880 5012
rect 252704 4972 252710 4984
rect 547874 4972 547880 4984
rect 547932 4972 547938 5024
rect 143534 4904 143540 4956
rect 143592 4944 143598 4956
rect 220998 4944 221004 4956
rect 143592 4916 221004 4944
rect 143592 4904 143598 4916
rect 220998 4904 221004 4916
rect 221056 4904 221062 4956
rect 229462 4904 229468 4956
rect 229520 4944 229526 4956
rect 241698 4944 241704 4956
rect 229520 4916 241704 4944
rect 229520 4904 229526 4916
rect 241698 4904 241704 4916
rect 241756 4904 241762 4956
rect 252554 4904 252560 4956
rect 252612 4944 252618 4956
rect 551462 4944 551468 4956
rect 252612 4916 551468 4944
rect 252612 4904 252618 4916
rect 551462 4904 551468 4916
rect 551520 4904 551526 4956
rect 132954 4836 132960 4888
rect 133012 4876 133018 4888
rect 219710 4876 219716 4888
rect 133012 4848 219716 4876
rect 133012 4836 133018 4848
rect 219710 4836 219716 4848
rect 219768 4836 219774 4888
rect 229646 4836 229652 4888
rect 229704 4876 229710 4888
rect 251174 4876 251180 4888
rect 229704 4848 251180 4876
rect 229704 4836 229710 4848
rect 251174 4836 251180 4848
rect 251232 4836 251238 4888
rect 252738 4836 252744 4888
rect 252796 4876 252802 4888
rect 554958 4876 554964 4888
rect 252796 4848 554964 4876
rect 252796 4836 252802 4848
rect 554958 4836 554964 4848
rect 555016 4836 555022 4888
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 203518 4808 203524 4820
rect 19484 4780 203524 4808
rect 19484 4768 19490 4780
rect 203518 4768 203524 4780
rect 203576 4768 203582 4820
rect 205082 4768 205088 4820
rect 205140 4808 205146 4820
rect 225138 4808 225144 4820
rect 205140 4780 225144 4808
rect 205140 4768 205146 4780
rect 225138 4768 225144 4780
rect 225196 4768 225202 4820
rect 229554 4768 229560 4820
rect 229612 4808 229618 4820
rect 252370 4808 252376 4820
rect 229612 4780 252376 4808
rect 229612 4768 229618 4780
rect 252370 4768 252376 4780
rect 252428 4768 252434 4820
rect 254946 4768 254952 4820
rect 255004 4808 255010 4820
rect 560846 4808 560852 4820
rect 255004 4780 560852 4808
rect 255004 4768 255010 4780
rect 560846 4768 560852 4780
rect 560904 4768 560910 4820
rect 228082 4088 228088 4140
rect 228140 4128 228146 4140
rect 229830 4128 229836 4140
rect 228140 4100 229836 4128
rect 228140 4088 228146 4100
rect 229830 4088 229836 4100
rect 229888 4088 229894 4140
rect 230566 4088 230572 4140
rect 230624 4128 230630 4140
rect 239398 4128 239404 4140
rect 230624 4100 239404 4128
rect 230624 4088 230630 4100
rect 239398 4088 239404 4100
rect 239456 4088 239462 4140
rect 242158 4088 242164 4140
rect 242216 4128 242222 4140
rect 259454 4128 259460 4140
rect 242216 4100 259460 4128
rect 242216 4088 242222 4100
rect 259454 4088 259460 4100
rect 259512 4088 259518 4140
rect 217962 4020 217968 4072
rect 218020 4060 218026 4072
rect 223942 4060 223948 4072
rect 218020 4032 223948 4060
rect 218020 4020 218026 4032
rect 223942 4020 223948 4032
rect 224000 4020 224006 4072
rect 231762 4020 231768 4072
rect 231820 4060 231826 4072
rect 231820 4032 233556 4060
rect 231820 4020 231826 4032
rect 95142 3952 95148 4004
rect 95200 3992 95206 4004
rect 149698 3992 149704 4004
rect 95200 3964 149704 3992
rect 95200 3952 95206 3964
rect 149698 3952 149704 3964
rect 149756 3952 149762 4004
rect 219250 3952 219256 4004
rect 219308 3992 219314 4004
rect 222838 3992 222844 4004
rect 219308 3964 222844 3992
rect 219308 3952 219314 3964
rect 222838 3952 222844 3964
rect 222896 3952 222902 4004
rect 227898 3952 227904 4004
rect 227956 3992 227962 4004
rect 233418 3992 233424 4004
rect 227956 3964 233424 3992
rect 227956 3952 227962 3964
rect 233418 3952 233424 3964
rect 233476 3952 233482 4004
rect 233528 3992 233556 4032
rect 234890 4020 234896 4072
rect 234948 4060 234954 4072
rect 258258 4060 258264 4072
rect 234948 4032 258264 4060
rect 234948 4020 234954 4032
rect 258258 4020 258264 4032
rect 258316 4020 258322 4072
rect 260650 3992 260656 4004
rect 233528 3964 260656 3992
rect 260650 3952 260656 3964
rect 260708 3952 260714 4004
rect 115198 3884 115204 3936
rect 115256 3924 115262 3936
rect 171778 3924 171784 3936
rect 115256 3896 171784 3924
rect 115256 3884 115262 3896
rect 171778 3884 171784 3896
rect 171836 3884 171842 3936
rect 186130 3884 186136 3936
rect 186188 3924 186194 3936
rect 224310 3924 224316 3936
rect 186188 3896 224316 3924
rect 186188 3884 186194 3896
rect 224310 3884 224316 3896
rect 224368 3884 224374 3936
rect 227990 3884 227996 3936
rect 228048 3924 228054 3936
rect 235810 3924 235816 3936
rect 228048 3896 235816 3924
rect 228048 3884 228054 3896
rect 235810 3884 235816 3896
rect 235868 3884 235874 3936
rect 236086 3884 236092 3936
rect 236144 3924 236150 3936
rect 239306 3924 239312 3936
rect 236144 3896 239312 3924
rect 236144 3884 236150 3896
rect 239306 3884 239312 3896
rect 239364 3884 239370 3936
rect 239398 3884 239404 3936
rect 239456 3924 239462 3936
rect 271230 3924 271236 3936
rect 239456 3896 271236 3924
rect 239456 3884 239462 3896
rect 271230 3884 271236 3896
rect 271288 3884 271294 3936
rect 112806 3816 112812 3868
rect 112864 3856 112870 3868
rect 169018 3856 169024 3868
rect 112864 3828 169024 3856
rect 112864 3816 112870 3828
rect 169018 3816 169024 3828
rect 169076 3816 169082 3868
rect 184934 3816 184940 3868
rect 184992 3856 184998 3868
rect 209038 3856 209044 3868
rect 184992 3828 209044 3856
rect 184992 3816 184998 3828
rect 209038 3816 209044 3828
rect 209096 3816 209102 3868
rect 219342 3816 219348 3868
rect 219400 3856 219406 3868
rect 264146 3856 264152 3868
rect 219400 3828 264152 3856
rect 219400 3816 219406 3828
rect 264146 3816 264152 3828
rect 264204 3816 264210 3868
rect 284294 3816 284300 3868
rect 284352 3856 284358 3868
rect 285030 3856 285036 3868
rect 284352 3828 285036 3856
rect 284352 3816 284358 3828
rect 285030 3816 285036 3828
rect 285088 3816 285094 3868
rect 82078 3748 82084 3800
rect 82136 3788 82142 3800
rect 138658 3788 138664 3800
rect 82136 3760 138664 3788
rect 82136 3748 82142 3760
rect 138658 3748 138664 3760
rect 138716 3748 138722 3800
rect 151814 3748 151820 3800
rect 151872 3788 151878 3800
rect 153010 3788 153016 3800
rect 151872 3760 153016 3788
rect 151872 3748 151878 3760
rect 153010 3748 153016 3760
rect 153068 3748 153074 3800
rect 168374 3748 168380 3800
rect 168432 3788 168438 3800
rect 207750 3788 207756 3800
rect 168432 3760 207756 3788
rect 168432 3748 168438 3760
rect 207750 3748 207756 3760
rect 207808 3748 207814 3800
rect 215662 3748 215668 3800
rect 215720 3788 215726 3800
rect 225598 3788 225604 3800
rect 215720 3760 225604 3788
rect 215720 3748 215726 3760
rect 225598 3748 225604 3760
rect 225656 3748 225662 3800
rect 233326 3748 233332 3800
rect 233384 3788 233390 3800
rect 296070 3788 296076 3800
rect 233384 3760 296076 3788
rect 233384 3748 233390 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 118786 3680 118792 3732
rect 118844 3720 118850 3732
rect 185578 3720 185584 3732
rect 118844 3692 185584 3720
rect 118844 3680 118850 3692
rect 185578 3680 185584 3692
rect 185636 3680 185642 3732
rect 214466 3680 214472 3732
rect 214524 3720 214530 3732
rect 226518 3720 226524 3732
rect 214524 3692 226524 3720
rect 214524 3680 214530 3692
rect 226518 3680 226524 3692
rect 226576 3680 226582 3732
rect 234246 3680 234252 3732
rect 234304 3720 234310 3732
rect 299658 3720 299664 3732
rect 234304 3692 299664 3720
rect 234304 3680 234310 3692
rect 299658 3680 299664 3692
rect 299716 3680 299722 3732
rect 135346 3612 135352 3664
rect 135404 3652 135410 3664
rect 207658 3652 207664 3664
rect 135404 3624 207664 3652
rect 135404 3612 135410 3624
rect 207658 3612 207664 3624
rect 207716 3612 207722 3664
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 227438 3652 227444 3664
rect 213420 3624 227444 3652
rect 213420 3612 213426 3624
rect 227438 3612 227444 3624
rect 227496 3612 227502 3664
rect 229002 3612 229008 3664
rect 229060 3652 229066 3664
rect 237006 3652 237012 3664
rect 229060 3624 237012 3652
rect 229060 3612 229066 3624
rect 237006 3612 237012 3624
rect 237064 3612 237070 3664
rect 239490 3612 239496 3664
rect 239548 3652 239554 3664
rect 335078 3652 335084 3664
rect 239548 3624 335084 3652
rect 239548 3612 239554 3624
rect 335078 3612 335084 3624
rect 335136 3612 335142 3664
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 88242 3584 88248 3596
rect 12400 3556 88248 3584
rect 12400 3544 12406 3556
rect 88242 3544 88248 3556
rect 88300 3544 88306 3596
rect 88978 3544 88984 3596
rect 89036 3544 89042 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 219526 3584 219532 3596
rect 129424 3556 219532 3584
rect 129424 3544 129430 3556
rect 219526 3544 219532 3556
rect 219584 3544 219590 3596
rect 229370 3544 229376 3596
rect 229428 3584 229434 3596
rect 246390 3584 246396 3596
rect 229428 3556 234200 3584
rect 229428 3544 229434 3556
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 88996 3516 89024 3544
rect 13596 3488 89024 3516
rect 13596 3476 13602 3488
rect 118694 3476 118700 3528
rect 118752 3516 118758 3528
rect 119890 3516 119896 3528
rect 118752 3488 119896 3516
rect 118752 3476 118758 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 219618 3516 219624 3528
rect 127032 3488 219624 3516
rect 127032 3476 127038 3488
rect 219618 3476 219624 3488
rect 219676 3476 219682 3528
rect 231118 3476 231124 3528
rect 231176 3516 231182 3528
rect 232222 3516 232228 3528
rect 231176 3488 232228 3516
rect 231176 3476 231182 3488
rect 232222 3476 232228 3488
rect 232280 3476 232286 3528
rect 234172 3516 234200 3556
rect 239324 3556 246396 3584
rect 236546 3516 236552 3528
rect 234172 3488 236552 3516
rect 236546 3476 236552 3488
rect 236604 3476 236610 3528
rect 44174 3408 44180 3460
rect 44232 3448 44238 3460
rect 45094 3448 45100 3460
rect 44232 3420 45100 3448
rect 44232 3408 44238 3420
rect 45094 3408 45100 3420
rect 45152 3408 45158 3460
rect 52546 3408 52552 3460
rect 52604 3448 52610 3460
rect 52604 3420 161474 3448
rect 52604 3408 52610 3420
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136450 3380 136456 3392
rect 135312 3352 136456 3380
rect 135312 3340 135318 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 161446 3380 161474 3420
rect 176654 3408 176660 3460
rect 176712 3448 176718 3460
rect 177850 3448 177856 3460
rect 176712 3420 177856 3448
rect 176712 3408 176718 3420
rect 177850 3408 177856 3420
rect 177908 3408 177914 3460
rect 182542 3408 182548 3460
rect 182600 3448 182606 3460
rect 223666 3448 223672 3460
rect 182600 3420 223672 3448
rect 182600 3408 182606 3420
rect 223666 3408 223672 3420
rect 223724 3408 223730 3460
rect 229186 3408 229192 3460
rect 229244 3448 229250 3460
rect 239324 3448 239352 3556
rect 246390 3544 246396 3556
rect 246448 3544 246454 3596
rect 257338 3544 257344 3596
rect 257396 3584 257402 3596
rect 465166 3584 465172 3596
rect 257396 3556 465172 3584
rect 257396 3544 257402 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 473354 3544 473360 3596
rect 473412 3584 473418 3596
rect 474182 3584 474188 3596
rect 473412 3556 474188 3584
rect 473412 3544 473418 3556
rect 474182 3544 474188 3556
rect 474240 3544 474246 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482462 3584 482468 3596
rect 481692 3556 482468 3584
rect 481692 3544 481698 3556
rect 482462 3544 482468 3556
rect 482520 3544 482526 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 490742 3584 490748 3596
rect 489972 3556 490748 3584
rect 489972 3544 489978 3556
rect 490742 3544 490748 3556
rect 490800 3544 490806 3596
rect 239398 3476 239404 3528
rect 239456 3516 239462 3528
rect 247586 3516 247592 3528
rect 239456 3488 247592 3516
rect 239456 3476 239462 3488
rect 247586 3476 247592 3488
rect 247644 3476 247650 3528
rect 248414 3476 248420 3528
rect 248472 3516 248478 3528
rect 501782 3516 501788 3528
rect 248472 3488 501788 3516
rect 248472 3476 248478 3488
rect 501782 3476 501788 3488
rect 501840 3476 501846 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 581822 3516 581828 3528
rect 581052 3488 581828 3516
rect 581052 3476 581058 3488
rect 581822 3476 581828 3488
rect 581880 3476 581886 3528
rect 229244 3420 239352 3448
rect 229244 3408 229250 3420
rect 255958 3408 255964 3460
rect 256016 3448 256022 3460
rect 530118 3448 530124 3460
rect 256016 3420 530124 3448
rect 256016 3408 256022 3420
rect 530118 3408 530124 3420
rect 530176 3408 530182 3460
rect 178770 3380 178776 3392
rect 161446 3352 178776 3380
rect 178770 3340 178776 3352
rect 178828 3340 178834 3392
rect 201494 3340 201500 3392
rect 201552 3380 201558 3392
rect 202690 3380 202696 3392
rect 201552 3352 202696 3380
rect 201552 3340 201558 3352
rect 202690 3340 202696 3352
rect 202748 3340 202754 3392
rect 221550 3340 221556 3392
rect 221608 3380 221614 3392
rect 225690 3380 225696 3392
rect 221608 3352 225696 3380
rect 221608 3340 221614 3352
rect 225690 3340 225696 3352
rect 225748 3340 225754 3392
rect 230106 3340 230112 3392
rect 230164 3380 230170 3392
rect 244090 3380 244096 3392
rect 230164 3352 244096 3380
rect 230164 3340 230170 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 299566 3340 299572 3392
rect 299624 3380 299630 3392
rect 300762 3380 300768 3392
rect 299624 3352 300768 3380
rect 299624 3340 299630 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 456886 3340 456892 3392
rect 456944 3380 456950 3392
rect 458082 3380 458088 3392
rect 456944 3352 458088 3380
rect 456944 3340 456950 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 229278 3272 229284 3324
rect 229336 3312 229342 3324
rect 229336 3284 234614 3312
rect 229336 3272 229342 3284
rect 20622 3204 20628 3256
rect 20680 3244 20686 3256
rect 25498 3244 25504 3256
rect 20680 3216 25504 3244
rect 20680 3204 20686 3216
rect 25498 3204 25504 3216
rect 25556 3204 25562 3256
rect 234586 3244 234614 3284
rect 236546 3272 236552 3324
rect 236604 3312 236610 3324
rect 239398 3312 239404 3324
rect 236604 3284 239404 3312
rect 236604 3272 236610 3284
rect 239398 3272 239404 3284
rect 239456 3272 239462 3324
rect 240778 3272 240784 3324
rect 240836 3312 240842 3324
rect 240836 3284 241514 3312
rect 240836 3272 240842 3284
rect 241486 3244 241514 3284
rect 248782 3244 248788 3256
rect 234586 3216 234752 3244
rect 241486 3216 248788 3244
rect 232498 3068 232504 3120
rect 232556 3108 232562 3120
rect 234614 3108 234620 3120
rect 232556 3080 234620 3108
rect 232556 3068 232562 3080
rect 234614 3068 234620 3080
rect 234672 3068 234678 3120
rect 234724 3108 234752 3216
rect 248782 3204 248788 3216
rect 248840 3204 248846 3256
rect 236638 3136 236644 3188
rect 236696 3176 236702 3188
rect 242894 3176 242900 3188
rect 236696 3148 242900 3176
rect 236696 3136 236702 3148
rect 242894 3136 242900 3148
rect 242952 3136 242958 3188
rect 249978 3108 249984 3120
rect 234724 3080 249984 3108
rect 249978 3068 249984 3080
rect 250036 3068 250042 3120
rect 227622 2864 227628 2916
rect 227680 2904 227686 2916
rect 231026 2904 231032 2916
rect 227680 2876 231032 2904
rect 227680 2864 227686 2876
rect 231026 2864 231032 2876
rect 231084 2864 231090 2916
rect 423674 1368 423680 1420
rect 423732 1408 423738 1420
rect 424962 1408 424968 1420
rect 423732 1380 424968 1408
rect 423732 1368 423738 1380
rect 424962 1368 424968 1380
rect 425020 1368 425026 1420
rect 448514 1368 448520 1420
rect 448572 1408 448578 1420
rect 449802 1408 449808 1420
rect 448572 1380 449808 1408
rect 448572 1368 448578 1380
rect 449802 1368 449808 1380
rect 449860 1368 449866 1420
rect 365714 1096 365720 1148
rect 365772 1136 365778 1148
rect 367002 1136 367008 1148
rect 365772 1108 367008 1136
rect 365772 1096 365778 1108
rect 367002 1096 367008 1108
rect 367060 1096 367066 1148
rect 390554 1096 390560 1148
rect 390612 1136 390618 1148
rect 391842 1136 391848 1148
rect 390612 1108 391848 1136
rect 390612 1096 390618 1108
rect 391842 1096 391848 1108
rect 391900 1096 391906 1148
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 405004 700544 405056 700596
rect 413652 700544 413704 700596
rect 154120 700476 154172 700528
rect 182824 700476 182876 700528
rect 296076 700476 296128 700528
rect 300124 700476 300176 700528
rect 409144 700476 409196 700528
rect 429844 700476 429896 700528
rect 137836 700408 137888 700460
rect 178684 700408 178736 700460
rect 188896 700408 188948 700460
rect 202788 700408 202840 700460
rect 293224 700408 293276 700460
rect 332508 700408 332560 700460
rect 403624 700408 403676 700460
rect 462320 700408 462372 700460
rect 105452 700340 105504 700392
rect 174544 700340 174596 700392
rect 188988 700340 189040 700392
rect 218980 700340 219032 700392
rect 291844 700340 291896 700392
rect 348792 700340 348844 700392
rect 399484 700340 399536 700392
rect 478512 700340 478564 700392
rect 89168 700272 89220 700324
rect 184204 700272 184256 700324
rect 188804 700272 188856 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 283012 700272 283064 700324
rect 295984 700272 296036 700324
rect 364984 700272 365036 700324
rect 406384 700272 406436 700324
rect 494796 700272 494848 700324
rect 509884 700272 509936 700324
rect 559656 700272 559708 700324
rect 170312 699660 170364 699712
rect 171784 699660 171836 699712
rect 395344 699660 395396 699712
rect 397460 699660 397512 699712
rect 286324 696940 286376 696992
rect 580172 696940 580224 696992
rect 508504 670692 508556 670744
rect 580172 670692 580224 670744
rect 512644 643084 512696 643136
rect 580172 643084 580224 643136
rect 501604 630640 501656 630692
rect 579988 630640 580040 630692
rect 504364 616836 504416 616888
rect 580172 616836 580224 616888
rect 297364 600108 297416 600160
rect 297916 600108 297968 600160
rect 78128 599972 78180 600024
rect 187240 599972 187292 600024
rect 408132 599972 408184 600024
rect 78036 599904 78088 599956
rect 187148 599904 187200 599956
rect 78588 599836 78640 599888
rect 187332 599836 187384 599888
rect 78220 599768 78272 599820
rect 186872 599768 186924 599820
rect 78496 599700 78548 599752
rect 186964 599700 187016 599752
rect 78404 599632 78456 599684
rect 187056 599632 187108 599684
rect 297456 598884 297508 598936
rect 408224 598884 408276 598936
rect 298008 598816 298060 598868
rect 407948 598816 408000 598868
rect 297548 598748 297600 598800
rect 407580 598748 407632 598800
rect 297272 598544 297324 598596
rect 298008 598544 298060 598596
rect 280988 597320 281040 597372
rect 335360 597320 335412 597372
rect 102876 597252 102928 597304
rect 212356 597252 212408 597304
rect 319996 597252 320048 597304
rect 427820 597252 427872 597304
rect 104808 597184 104860 597236
rect 214840 597184 214892 597236
rect 326160 597184 326212 597236
rect 434720 597184 434772 597236
rect 100668 597116 100720 597168
rect 209964 597116 210016 597168
rect 211068 597116 211120 597168
rect 318708 597116 318760 597168
rect 426440 597116 426492 597168
rect 99288 597048 99340 597100
rect 208952 597048 209004 597100
rect 324412 597048 324464 597100
rect 434720 597048 434772 597100
rect 102048 596980 102100 597032
rect 211160 596980 211212 597032
rect 212448 596980 212500 597032
rect 213828 596980 213880 597032
rect 284576 596980 284628 597032
rect 322940 596980 322992 597032
rect 433340 596980 433392 597032
rect 106188 596912 106240 596964
rect 215760 596912 215812 596964
rect 284392 596912 284444 596964
rect 320916 596912 320968 596964
rect 430580 596912 430632 596964
rect 103428 596844 103480 596896
rect 213828 596844 213880 596896
rect 214840 596844 214892 596896
rect 284484 596844 284536 596896
rect 299296 596844 299348 596896
rect 313280 596844 313332 596896
rect 97908 596776 97960 596828
rect 207848 596776 207900 596828
rect 212448 596776 212500 596828
rect 283196 596776 283248 596828
rect 299204 596776 299256 596828
rect 314660 596776 314712 596828
rect 281080 596708 281132 596760
rect 317696 596708 317748 596760
rect 318708 596708 318760 596760
rect 283104 596640 283156 596692
rect 320088 596640 320140 596692
rect 429200 596844 429252 596896
rect 283196 596572 283248 596624
rect 320916 596572 320968 596624
rect 140688 596504 140740 596556
rect 172152 596504 172204 596556
rect 284300 596504 284352 596556
rect 322204 596504 322256 596556
rect 431960 596776 432012 596828
rect 407948 596504 408000 596556
rect 422576 596504 422628 596556
rect 136548 596436 136600 596488
rect 173348 596436 173400 596488
rect 281540 596436 281592 596488
rect 319996 596436 320048 596488
rect 408132 596436 408184 596488
rect 423680 596436 423732 596488
rect 131028 596368 131080 596420
rect 171876 596368 171928 596420
rect 212356 596368 212408 596420
rect 284300 596368 284352 596420
rect 284576 596368 284628 596420
rect 322940 596368 322992 596420
rect 408224 596368 408276 596420
rect 425060 596368 425112 596420
rect 79784 596300 79836 596352
rect 92480 596300 92532 596352
rect 126888 596300 126940 596352
rect 173256 596300 173308 596352
rect 188620 596300 188672 596352
rect 202880 596300 202932 596352
rect 208952 596300 209004 596352
rect 281540 596300 281592 596352
rect 284484 596300 284536 596352
rect 324412 596300 324464 596352
rect 406476 596300 406528 596352
rect 434720 596300 434772 596352
rect 79968 596232 80020 596284
rect 94044 596232 94096 596284
rect 121368 596232 121420 596284
rect 171968 596232 172020 596284
rect 188712 596232 188764 596284
rect 204352 596232 204404 596284
rect 211068 596232 211120 596284
rect 283104 596232 283156 596284
rect 284392 596232 284444 596284
rect 326160 596232 326212 596284
rect 409420 596232 409472 596284
rect 444380 596232 444432 596284
rect 79876 596164 79928 596216
rect 95240 596164 95292 596216
rect 115848 596164 115900 596216
rect 172060 596164 172112 596216
rect 188528 596164 188580 596216
rect 204260 596164 204312 596216
rect 207848 596164 207900 596216
rect 281080 596164 281132 596216
rect 299388 596164 299440 596216
rect 311900 596164 311952 596216
rect 409236 596164 409288 596216
rect 455420 596164 455472 596216
rect 282184 592628 282236 592680
rect 440240 592628 440292 592680
rect 285036 590656 285088 590708
rect 580172 590656 580224 590708
rect 289084 589908 289136 589960
rect 329840 589908 329892 589960
rect 284944 588548 284996 588600
rect 339500 588548 339552 588600
rect 287704 587188 287756 587240
rect 324320 587188 324372 587240
rect 282276 587120 282328 587172
rect 449900 587120 449952 587172
rect 286416 585828 286468 585880
rect 360200 585828 360252 585880
rect 297180 585760 297232 585812
rect 407672 585760 407724 585812
rect 78312 584400 78364 584452
rect 186780 584400 186832 584452
rect 298744 584400 298796 584452
rect 354680 584400 354732 584452
rect 291936 582972 291988 583024
rect 349160 582972 349212 583024
rect 111708 581612 111760 581664
rect 188344 581612 188396 581664
rect 226248 581612 226300 581664
rect 281632 581612 281684 581664
rect 289176 581612 289228 581664
rect 345020 581612 345072 581664
rect 251088 580524 251140 580576
rect 281724 580524 281776 580576
rect 245568 580456 245620 580508
rect 281816 580456 281868 580508
rect 241428 580388 241480 580440
rect 282092 580388 282144 580440
rect 190000 580320 190052 580372
rect 215300 580320 215352 580372
rect 235908 580320 235960 580372
rect 281908 580320 281960 580372
rect 189908 580252 189960 580304
rect 219440 580252 219492 580304
rect 231768 580252 231820 580304
rect 282000 580252 282052 580304
rect 282368 580252 282420 580304
rect 459560 580252 459612 580304
rect 516784 576852 516836 576904
rect 580172 576852 580224 576904
rect 3332 565836 3384 565888
rect 32404 565836 32456 565888
rect 507124 563048 507176 563100
rect 580172 563048 580224 563100
rect 3148 553392 3200 553444
rect 22744 553392 22796 553444
rect 511264 536800 511316 536852
rect 579896 536800 579948 536852
rect 3332 527144 3384 527196
rect 14464 527144 14516 527196
rect 293868 526736 293920 526788
rect 297272 526736 297324 526788
rect 298008 526736 298060 526788
rect 187332 525784 187384 525836
rect 187700 525784 187752 525836
rect 514024 524424 514076 524476
rect 580172 524424 580224 524476
rect 502984 510620 503036 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 10324 500964 10376 501016
rect 287796 498788 287848 498840
rect 296996 498788 297048 498840
rect 297824 498788 297876 498840
rect 187056 493348 187108 493400
rect 186688 493212 186740 493264
rect 187056 493212 187108 493264
rect 186872 493076 186924 493128
rect 78496 489812 78548 489864
rect 187700 489812 187752 489864
rect 297456 489812 297508 489864
rect 297732 489812 297784 489864
rect 407672 489812 407724 489864
rect 77668 489744 77720 489796
rect 187240 489744 187292 489796
rect 78404 489676 78456 489728
rect 187056 489676 187108 489728
rect 78312 489608 78364 489660
rect 187332 489608 187384 489660
rect 78128 489540 78180 489592
rect 186964 489540 187016 489592
rect 77760 489472 77812 489524
rect 186780 489472 186832 489524
rect 78036 489404 78088 489456
rect 186872 489404 186924 489456
rect 78588 489336 78640 489388
rect 187148 489336 187200 489388
rect 173348 489200 173400 489252
rect 253664 489200 253716 489252
rect 218060 489132 218112 489184
rect 405004 489132 405056 489184
rect 186872 488724 186924 488776
rect 187608 488724 187660 488776
rect 187240 488656 187292 488708
rect 187516 488656 187568 488708
rect 187056 488588 187108 488640
rect 187424 488588 187476 488640
rect 186780 488520 186832 488572
rect 187240 488520 187292 488572
rect 79784 488452 79836 488504
rect 92940 488452 92992 488504
rect 188620 488452 188672 488504
rect 297088 488452 297140 488504
rect 297548 488452 297600 488504
rect 297732 488452 297784 488504
rect 298008 488452 298060 488504
rect 408224 488452 408276 488504
rect 425060 488452 425112 488504
rect 79968 488384 80020 488436
rect 94228 488384 94280 488436
rect 188528 488384 188580 488436
rect 204720 488384 204772 488436
rect 292028 488384 292080 488436
rect 297640 488384 297692 488436
rect 407856 488384 407908 488436
rect 408132 488384 408184 488436
rect 423680 488384 423732 488436
rect 79876 488316 79928 488368
rect 95332 488316 95384 488368
rect 298008 488316 298060 488368
rect 407764 488316 407816 488368
rect 407948 488316 408000 488368
rect 422576 488316 422628 488368
rect 298100 488248 298152 488300
rect 299296 488248 299348 488300
rect 314292 488248 314344 488300
rect 408132 488248 408184 488300
rect 188620 488180 188672 488232
rect 202880 488180 202932 488232
rect 188712 488112 188764 488164
rect 204904 488112 204956 488164
rect 188804 488044 188856 488096
rect 220084 488044 220136 488096
rect 105728 487976 105780 488028
rect 215760 487976 215812 488028
rect 230572 487976 230624 488028
rect 287796 487976 287848 488028
rect 104808 487908 104860 487960
rect 214840 487908 214892 487960
rect 219808 487908 219860 487960
rect 283012 487908 283064 487960
rect 103428 487840 103480 487892
rect 213736 487840 213788 487892
rect 232596 487840 232648 487892
rect 299204 488180 299256 488232
rect 315396 488180 315448 488232
rect 408224 488180 408276 488232
rect 297548 488112 297600 488164
rect 408316 488112 408368 488164
rect 101128 487772 101180 487824
rect 211160 487772 211212 487824
rect 212448 487772 212500 487824
rect 232504 487772 232556 487824
rect 298100 487772 298152 487824
rect 312544 487772 312596 487824
rect 313004 487772 313056 487824
rect 407948 487772 408000 487824
rect 326620 487636 326672 487688
rect 434720 487636 434772 487688
rect 319444 487568 319496 487620
rect 427820 487568 427872 487620
rect 318064 487500 318116 487552
rect 426440 487500 426492 487552
rect 97816 487432 97868 487484
rect 207664 487432 207716 487484
rect 214840 487432 214892 487484
rect 228364 487432 228416 487484
rect 319996 487432 320048 487484
rect 429200 487432 429252 487484
rect 102416 487364 102468 487416
rect 212356 487364 212408 487416
rect 212448 487364 212500 487416
rect 226984 487364 227036 487416
rect 322940 487364 322992 487416
rect 433340 487364 433392 487416
rect 98920 487296 98972 487348
rect 208860 487296 208912 487348
rect 213736 487296 213788 487348
rect 229744 487296 229796 487348
rect 324412 487296 324464 487348
rect 434720 487296 434772 487348
rect 204720 487228 204772 487280
rect 222844 487228 222896 487280
rect 322204 487228 322256 487280
rect 432144 487228 432196 487280
rect 100024 487160 100076 487212
rect 210424 487160 210476 487212
rect 215760 487160 215812 487212
rect 244280 487160 244332 487212
rect 320824 487160 320876 487212
rect 430580 487160 430632 487212
rect 436744 487160 436796 487212
rect 465080 487160 465132 487212
rect 299388 487092 299440 487144
rect 311900 487092 311952 487144
rect 312544 487092 312596 487144
rect 246488 486616 246540 486668
rect 249800 486616 249852 486668
rect 208860 486548 208912 486600
rect 238024 486548 238076 486600
rect 244924 486548 244976 486600
rect 324412 486548 324464 486600
rect 187700 486480 187752 486532
rect 235264 486480 235316 486532
rect 248420 486480 248472 486532
rect 409420 486480 409472 486532
rect 216772 486412 216824 486464
rect 542360 486412 542412 486464
rect 243820 485800 243872 485852
rect 244648 485800 244700 485852
rect 239404 485188 239456 485240
rect 319996 485188 320048 485240
rect 172152 485120 172204 485172
rect 254952 485120 255004 485172
rect 253940 485052 253992 485104
rect 409328 485052 409380 485104
rect 221464 484372 221516 484424
rect 580172 484372 580224 484424
rect 244280 484304 244332 484356
rect 326620 484304 326672 484356
rect 212356 483692 212408 483744
rect 242164 483692 242216 483744
rect 251180 483692 251232 483744
rect 409236 483692 409288 483744
rect 216956 483624 217008 483676
rect 580264 483624 580316 483676
rect 105820 482332 105872 482384
rect 234620 482332 234672 482384
rect 236092 482332 236144 482384
rect 434720 482332 434772 482384
rect 216680 482264 216732 482316
rect 501604 482264 501656 482316
rect 173256 481108 173308 481160
rect 250812 481108 250864 481160
rect 243544 481040 243596 481092
rect 322940 481040 322992 481092
rect 247868 480972 247920 481024
rect 360200 480972 360252 481024
rect 215300 480904 215352 480956
rect 516784 480904 516836 480956
rect 126888 479680 126940 479732
rect 240876 479680 240928 479732
rect 238852 479612 238904 479664
rect 339500 479612 339552 479664
rect 240784 479544 240836 479596
rect 320824 479544 320876 479596
rect 215484 479476 215536 479528
rect 514024 479476 514076 479528
rect 241428 478932 241480 478984
rect 242256 478932 242308 478984
rect 172060 478252 172112 478304
rect 248512 478252 248564 478304
rect 246580 478184 246632 478236
rect 354680 478184 354732 478236
rect 218244 478116 218296 478168
rect 395344 478116 395396 478168
rect 235264 477436 235316 477488
rect 293316 477436 293368 477488
rect 218152 476824 218204 476876
rect 403624 476824 403676 476876
rect 220728 476756 220780 476808
rect 229836 476756 229888 476808
rect 243636 476756 243688 476808
rect 459560 476756 459612 476808
rect 234804 476076 234856 476128
rect 235264 476076 235316 476128
rect 236552 475464 236604 475516
rect 318064 475464 318116 475516
rect 77944 475396 77996 475448
rect 229928 475396 229980 475448
rect 236276 475396 236328 475448
rect 329840 475396 329892 475448
rect 217140 475328 217192 475380
rect 527180 475328 527232 475380
rect 3240 474716 3292 474768
rect 40684 474716 40736 474768
rect 241612 474648 241664 474700
rect 242164 474648 242216 474700
rect 322204 474648 322256 474700
rect 173164 474104 173216 474156
rect 245660 474104 245712 474156
rect 237748 474036 237800 474088
rect 335360 474036 335412 474088
rect 215668 473968 215720 474020
rect 512644 473968 512696 474020
rect 237564 473288 237616 473340
rect 238024 473288 238076 473340
rect 319444 473288 319496 473340
rect 235908 473016 235960 473068
rect 240968 473016 241020 473068
rect 216588 472744 216640 472796
rect 235540 472744 235592 472796
rect 32404 472676 32456 472728
rect 224316 472676 224368 472728
rect 236000 472676 236052 472728
rect 324320 472676 324372 472728
rect 215392 472608 215444 472660
rect 511264 472608 511316 472660
rect 40684 471248 40736 471300
rect 224500 471248 224552 471300
rect 237472 471248 237524 471300
rect 440240 471248 440292 471300
rect 214012 470568 214064 470620
rect 579988 470568 580040 470620
rect 10324 469888 10376 469940
rect 224684 469888 224736 469940
rect 240324 469888 240376 469940
rect 455420 469888 455472 469940
rect 217324 469820 217376 469872
rect 509884 469820 509936 469872
rect 219624 468596 219676 468648
rect 296076 468596 296128 468648
rect 218336 468528 218388 468580
rect 399484 468528 399536 468580
rect 22744 468460 22796 468512
rect 223764 468460 223816 468512
rect 239036 468460 239088 468512
rect 449900 468460 449952 468512
rect 178684 467236 178736 467288
rect 221372 467236 221424 467288
rect 218428 467168 218480 467220
rect 409144 467168 409196 467220
rect 121368 467100 121420 467152
rect 239496 467100 239548 467152
rect 244556 467100 244608 467152
rect 470600 467100 470652 467152
rect 136548 465808 136600 465860
rect 243360 465808 243412 465860
rect 217508 465740 217560 465792
rect 406384 465740 406436 465792
rect 243084 465672 243136 465724
rect 436744 465672 436796 465724
rect 231492 464448 231544 464500
rect 311900 464448 311952 464500
rect 4068 464380 4120 464432
rect 224224 464380 224276 464432
rect 239220 464380 239272 464432
rect 444380 464380 444432 464432
rect 215852 464312 215904 464364
rect 504364 464312 504416 464364
rect 219716 463156 219768 463208
rect 282920 463156 282972 463208
rect 240508 463088 240560 463140
rect 345020 463088 345072 463140
rect 230756 463020 230808 463072
rect 408040 463020 408092 463072
rect 216864 462952 216916 463004
rect 508504 462952 508556 463004
rect 2872 462340 2924 462392
rect 225604 462340 225656 462392
rect 219900 461796 219952 461848
rect 291844 461796 291896 461848
rect 131028 461728 131080 461780
rect 242072 461728 242124 461780
rect 71780 461660 71832 461712
rect 221556 461660 221608 461712
rect 241796 461660 241848 461712
rect 349160 461660 349212 461712
rect 215760 461592 215812 461644
rect 507124 461592 507176 461644
rect 207664 460844 207716 460896
rect 236552 460844 236604 460896
rect 218612 460300 218664 460352
rect 293224 460300 293276 460352
rect 14464 460232 14516 460284
rect 224040 460232 224092 460284
rect 245844 460232 245896 460284
rect 406476 460232 406528 460284
rect 214196 460164 214248 460216
rect 502984 460164 503036 460216
rect 210424 459484 210476 459536
rect 239128 459484 239180 459536
rect 239404 459484 239456 459536
rect 203524 459416 203576 459468
rect 231584 459416 231636 459468
rect 299664 458940 299716 458992
rect 321284 458940 321336 458992
rect 171968 458872 172020 458924
rect 249800 458872 249852 458924
rect 251824 458872 251876 458924
rect 371516 458872 371568 458924
rect 40040 458804 40092 458856
rect 221004 458804 221056 458856
rect 247040 458804 247092 458856
rect 379888 458804 379940 458856
rect 299388 458736 299440 458788
rect 329656 458736 329708 458788
rect 299480 458668 299532 458720
rect 342536 458668 342588 458720
rect 296076 458600 296128 458652
rect 346400 458600 346452 458652
rect 299572 458532 299624 458584
rect 350908 458532 350960 458584
rect 298928 458464 298980 458516
rect 359280 458464 359332 458516
rect 298008 458396 298060 458448
rect 367652 458396 367704 458448
rect 246304 458328 246356 458380
rect 363144 458328 363196 458380
rect 293316 458260 293368 458312
rect 309048 458260 309100 458312
rect 355968 458192 356020 458244
rect 376024 458192 376076 458244
rect 174544 457512 174596 457564
rect 220820 457512 220872 457564
rect 6920 457444 6972 457496
rect 222016 457444 222068 457496
rect 227352 457444 227404 457496
rect 355968 457444 356020 457496
rect 222936 457240 222988 457292
rect 317420 457240 317472 457292
rect 228456 457172 228508 457224
rect 325792 457172 325844 457224
rect 236368 457104 236420 457156
rect 338028 457104 338080 457156
rect 228548 457036 228600 457088
rect 334164 457036 334216 457088
rect 247132 456968 247184 457020
rect 354772 456968 354824 457020
rect 223028 456900 223080 456952
rect 383752 456900 383804 456952
rect 223856 456764 223908 456816
rect 224316 456764 224368 456816
rect 385316 456832 385368 456884
rect 299020 456764 299072 456816
rect 580172 456764 580224 456816
rect 299756 456016 299808 456068
rect 300768 456016 300820 456068
rect 235080 455948 235132 456000
rect 312636 455948 312688 456000
rect 252744 455880 252796 455932
rect 385132 455880 385184 455932
rect 251916 455812 251968 455864
rect 385224 455812 385276 455864
rect 250536 455744 250588 455796
rect 384120 455744 384172 455796
rect 244464 455676 244516 455728
rect 384212 455676 384264 455728
rect 298836 455608 298888 455660
rect 300308 455608 300360 455660
rect 300768 455608 300820 455660
rect 385040 455608 385092 455660
rect 237748 455540 237800 455592
rect 384028 455540 384080 455592
rect 214288 455472 214340 455524
rect 384304 455472 384356 455524
rect 214472 455404 214524 455456
rect 580264 455404 580316 455456
rect 299848 455336 299900 455388
rect 304172 455336 304224 455388
rect 249248 454860 249300 454912
rect 299848 454860 299900 454912
rect 235356 454792 235408 454844
rect 299572 454792 299624 454844
rect 235264 454724 235316 454776
rect 299480 454724 299532 454776
rect 219072 454656 219124 454708
rect 295984 454656 296036 454708
rect 182824 453432 182876 453484
rect 221740 453432 221792 453484
rect 215944 453364 215996 453416
rect 285036 453364 285088 453416
rect 214656 453296 214708 453348
rect 299020 453296 299072 453348
rect 237564 452548 237616 452600
rect 237840 452548 237892 452600
rect 243176 452344 243228 452396
rect 247040 452344 247092 452396
rect 219716 452276 219768 452328
rect 219992 452276 220044 452328
rect 255872 452276 255924 452328
rect 284392 452276 284444 452328
rect 254584 452208 254636 452260
rect 284484 452208 284536 452260
rect 253296 452140 253348 452192
rect 284576 452140 284628 452192
rect 247316 452072 247368 452124
rect 281540 452072 281592 452124
rect 246028 452004 246080 452056
rect 281080 452004 281132 452056
rect 171784 451936 171836 451988
rect 220728 451936 220780 451988
rect 234620 451936 234672 451988
rect 235632 451936 235684 451988
rect 239036 451936 239088 451988
rect 240048 451936 240100 451988
rect 240324 451936 240376 451988
rect 241336 451936 241388 451988
rect 247776 451936 247828 451988
rect 299388 451936 299440 451988
rect 217324 451868 217376 451920
rect 286324 451868 286376 451920
rect 214840 451256 214892 451308
rect 221464 451256 221516 451308
rect 233976 451256 234028 451308
rect 297640 451256 297692 451308
rect 228364 451188 228416 451240
rect 244280 451188 244332 451240
rect 189080 450916 189132 450968
rect 230848 450916 230900 450968
rect 188436 450848 188488 450900
rect 234252 450848 234304 450900
rect 187516 450780 187568 450832
rect 233424 450780 233476 450832
rect 256056 450780 256108 450832
rect 293316 450780 293368 450832
rect 187240 450712 187292 450764
rect 233792 450712 233844 450764
rect 254768 450712 254820 450764
rect 298008 450712 298060 450764
rect 187332 450644 187384 450696
rect 234068 450644 234120 450696
rect 244280 450644 244332 450696
rect 244924 450644 244976 450696
rect 255688 450644 255740 450696
rect 299756 450644 299808 450696
rect 187424 450576 187476 450628
rect 255412 450576 255464 450628
rect 187608 450508 187660 450560
rect 255320 450508 255372 450560
rect 230112 449896 230164 449948
rect 293224 449896 293276 449948
rect 3516 449828 3568 449880
rect 223028 449828 223080 449880
rect 234252 449828 234304 449880
rect 234528 449828 234580 449880
rect 297180 449828 297232 449880
rect 229744 449760 229796 449812
rect 242992 449760 243044 449812
rect 243544 449760 243596 449812
rect 253848 449760 253900 449812
rect 281816 449760 281868 449812
rect 187148 449692 187200 449744
rect 232688 449692 232740 449744
rect 252560 449692 252612 449744
rect 282092 449692 282144 449744
rect 189908 449624 189960 449676
rect 247408 449624 247460 449676
rect 251272 449624 251324 449676
rect 281908 449624 281960 449676
rect 190000 449556 190052 449608
rect 246120 449556 246172 449608
rect 249984 449556 250036 449608
rect 282000 449556 282052 449608
rect 188344 449488 188396 449540
rect 247224 449488 247276 449540
rect 250720 449488 250772 449540
rect 283196 449488 283248 449540
rect 252008 449420 252060 449472
rect 284300 449420 284352 449472
rect 140688 449352 140740 449404
rect 244648 449352 244700 449404
rect 248696 449352 248748 449404
rect 281632 449352 281684 449404
rect 115848 449284 115900 449336
rect 238208 449284 238260 449336
rect 249432 449284 249484 449336
rect 283104 449284 283156 449336
rect 111708 449216 111760 449268
rect 236920 449216 236972 449268
rect 246764 449216 246816 449268
rect 298928 449216 298980 449268
rect 3884 449148 3936 449200
rect 223120 449148 223172 449200
rect 241520 449148 241572 449200
rect 298836 449148 298888 449200
rect 204904 449080 204956 449132
rect 232596 449080 232648 449132
rect 255136 449080 255188 449132
rect 281724 449080 281776 449132
rect 186964 449012 187016 449064
rect 233056 449012 233108 449064
rect 171876 448944 171928 448996
rect 252376 448944 252428 448996
rect 252192 448604 252244 448656
rect 293316 448604 293368 448656
rect 222752 448536 222804 448588
rect 223028 448536 223080 448588
rect 247040 448536 247092 448588
rect 293408 448536 293460 448588
rect 23480 448468 23532 448520
rect 222200 448468 222252 448520
rect 222936 448468 222988 448520
rect 233056 448400 233108 448452
rect 297732 448468 297784 448520
rect 222844 448332 222896 448384
rect 231952 448332 232004 448384
rect 232504 448332 232556 448384
rect 232688 448332 232740 448384
rect 297364 448400 297416 448452
rect 240416 448332 240468 448384
rect 240784 448332 240836 448384
rect 233792 448264 233844 448316
rect 239404 448264 239456 448316
rect 184204 448196 184256 448248
rect 221648 448196 221700 448248
rect 226984 448196 227036 448248
rect 240416 448196 240468 448248
rect 3700 448128 3752 448180
rect 222936 448128 222988 448180
rect 233424 448128 233476 448180
rect 297824 448332 297876 448384
rect 297456 448264 297508 448316
rect 3976 448060 4028 448112
rect 223488 448060 223540 448112
rect 239404 448060 239456 448112
rect 255320 448196 255372 448248
rect 256240 448196 256292 448248
rect 297548 448196 297600 448248
rect 3424 447992 3476 448044
rect 222384 447992 222436 448044
rect 3608 447924 3660 447976
rect 222568 447924 222620 447976
rect 236736 447924 236788 447976
rect 251824 447924 251876 447976
rect 3792 447856 3844 447908
rect 223304 447856 223356 447908
rect 231768 447856 231820 447908
rect 239680 447856 239732 447908
rect 248880 447856 248932 447908
rect 280988 447856 281040 447908
rect 3240 447788 3292 447840
rect 224776 447788 224828 447840
rect 226248 447788 226300 447840
rect 238392 447788 238444 447840
rect 245660 447788 245712 447840
rect 296076 447788 296128 447840
rect 213184 447720 213236 447772
rect 219164 447720 219216 447772
rect 245844 447720 245896 447772
rect 246396 447720 246448 447772
rect 211712 447652 211764 447704
rect 218796 447652 218848 447704
rect 219440 447652 219492 447704
rect 219900 447652 219952 447704
rect 246028 447652 246080 447704
rect 246856 447652 246908 447704
rect 212816 447584 212868 447636
rect 212632 447516 212684 447568
rect 212264 447448 212316 447500
rect 214012 447312 214064 447364
rect 215024 447312 215076 447364
rect 215668 447312 215720 447364
rect 216496 447312 216548 447364
rect 214196 447244 214248 447296
rect 215208 447244 215260 447296
rect 215852 447244 215904 447296
rect 216312 447244 216364 447296
rect 215300 447176 215352 447228
rect 216128 447176 216180 447228
rect 217140 447312 217192 447364
rect 217600 447312 217652 447364
rect 218060 447312 218112 447364
rect 218888 447312 218940 447364
rect 241888 447584 241940 447636
rect 246304 447584 246356 447636
rect 221004 447516 221056 447568
rect 221832 447516 221884 447568
rect 240600 447516 240652 447568
rect 298008 447516 298060 447568
rect 296352 447448 296404 447500
rect 219164 447380 219216 447432
rect 296628 447380 296680 447432
rect 296444 447312 296496 447364
rect 218244 447244 218296 447296
rect 218704 447244 218756 447296
rect 218796 447244 218848 447296
rect 296168 447244 296220 447296
rect 296260 447176 296312 447228
rect 213736 447108 213788 447160
rect 299204 447108 299256 447160
rect 232044 447040 232096 447092
rect 232504 447040 232556 447092
rect 252928 447040 252980 447092
rect 282368 447040 282420 447092
rect 255320 446972 255372 447024
rect 286416 446972 286468 447024
rect 250352 446904 250404 446956
rect 282276 446904 282328 446956
rect 224960 446836 225012 446888
rect 225604 446836 225656 446888
rect 243728 446836 243780 446888
rect 246672 446836 246724 446888
rect 247776 446836 247828 446888
rect 282184 446836 282236 446888
rect 3700 446768 3752 446820
rect 227536 446768 227588 446820
rect 250168 446768 250220 446820
rect 284944 446768 284996 446820
rect 221648 446700 221700 446752
rect 248604 446700 248656 446752
rect 251456 446700 251508 446752
rect 289176 446700 289228 446752
rect 3424 446632 3476 446684
rect 228640 446632 228692 446684
rect 252744 446632 252796 446684
rect 291936 446632 291988 446684
rect 4988 446564 5040 446616
rect 225512 446564 225564 446616
rect 246304 446564 246356 446616
rect 287704 446564 287756 446616
rect 216588 446496 216640 446548
rect 227168 446496 227220 446548
rect 247592 446496 247644 446548
rect 289084 446496 289136 446548
rect 188896 446428 188948 446480
rect 220360 446428 220412 446480
rect 238944 446428 238996 446480
rect 243636 446428 243688 446480
rect 244832 446428 244884 446480
rect 252652 446428 252704 446480
rect 256608 446428 256660 446480
rect 299848 446428 299900 446480
rect 188988 446360 189040 446412
rect 220544 446360 220596 446412
rect 229928 446360 229980 446412
rect 230664 446360 230716 446412
rect 233240 446360 233292 446412
rect 251916 446360 251968 446412
rect 254032 446360 254084 446412
rect 298744 446360 298796 446412
rect 212080 446292 212132 446344
rect 299020 446292 299072 446344
rect 213368 446224 213420 446276
rect 296536 446224 296588 446276
rect 214104 446156 214156 446208
rect 298560 446156 298612 446208
rect 4896 446088 4948 446140
rect 226064 446088 226116 446140
rect 234344 446088 234396 446140
rect 255596 446088 255648 446140
rect 3884 446020 3936 446072
rect 226984 446020 227036 446072
rect 231400 446020 231452 446072
rect 255412 446020 255464 446072
rect 224960 445952 225012 446004
rect 254308 445952 254360 446004
rect 4804 445884 4856 445936
rect 228824 445884 228876 445936
rect 239312 445884 239364 445936
rect 3792 445816 3844 445868
rect 227720 445816 227772 445868
rect 229836 445816 229888 445868
rect 237104 445816 237156 445868
rect 242624 445816 242676 445868
rect 243452 445816 243504 445868
rect 243636 445884 243688 445936
rect 244832 445884 244884 445936
rect 249892 445884 249944 445936
rect 245016 445816 245068 445868
rect 248052 445816 248104 445868
rect 219348 445748 219400 445800
rect 225144 445748 225196 445800
rect 232872 445748 232924 445800
rect 227904 445680 227956 445732
rect 228456 445680 228508 445732
rect 244832 445748 244884 445800
rect 246580 445748 246632 445800
rect 245660 445680 245712 445732
rect 211528 445340 211580 445392
rect 220084 445340 220136 445392
rect 221096 445340 221148 445392
rect 221740 445340 221792 445392
rect 247132 445340 247184 445392
rect 248328 445340 248380 445392
rect 196716 445272 196768 445324
rect 226800 445272 226852 445324
rect 98644 445204 98696 445256
rect 225696 445204 225748 445256
rect 229560 445272 229612 445324
rect 267004 445272 267056 445324
rect 265900 445204 265952 445256
rect 199568 445136 199620 445188
rect 226248 445136 226300 445188
rect 234712 445136 234764 445188
rect 235356 445136 235408 445188
rect 236276 445136 236328 445188
rect 237288 445136 237340 445188
rect 238760 445136 238812 445188
rect 239220 445136 239272 445188
rect 240508 445136 240560 445188
rect 241152 445136 241204 445188
rect 241796 445136 241848 445188
rect 242440 445136 242492 445188
rect 243084 445136 243136 445188
rect 243912 445136 243964 445188
rect 244372 445136 244424 445188
rect 245568 445136 245620 445188
rect 247316 445136 247368 445188
rect 248144 445136 248196 445188
rect 248420 445136 248472 445188
rect 249064 445136 249116 445188
rect 251824 445136 251876 445188
rect 293868 445136 293920 445188
rect 3976 445068 4028 445120
rect 216588 445068 216640 445120
rect 216772 445068 216824 445120
rect 217784 445068 217836 445120
rect 218612 445068 218664 445120
rect 219256 445068 219308 445120
rect 220820 445068 220872 445120
rect 221280 445068 221332 445120
rect 224224 445068 224276 445120
rect 224684 445068 224736 445120
rect 238852 445068 238904 445120
rect 239864 445068 239916 445120
rect 244096 445068 244148 445120
rect 293684 445068 293736 445120
rect 3240 445000 3292 445052
rect 219348 445000 219400 445052
rect 248604 445000 248656 445052
rect 299480 445000 299532 445052
rect 213000 444932 213052 444984
rect 265716 444932 265768 444984
rect 199476 444864 199528 444916
rect 227352 444864 227404 444916
rect 240232 444864 240284 444916
rect 293592 444864 293644 444916
rect 199384 444796 199436 444848
rect 228456 444796 228508 444848
rect 235448 444796 235500 444848
rect 293500 444796 293552 444848
rect 211896 444728 211948 444780
rect 269856 444728 269908 444780
rect 211344 444660 211396 444712
rect 217048 444592 217100 444644
rect 217324 444592 217376 444644
rect 220084 444660 220136 444712
rect 271236 444660 271288 444712
rect 196624 444524 196676 444576
rect 273996 444592 274048 444644
rect 227904 444524 227956 444576
rect 230480 444524 230532 444576
rect 298652 444524 298704 444576
rect 213920 444456 213972 444508
rect 295892 444456 295944 444508
rect 200856 444388 200908 444440
rect 229008 444388 229060 444440
rect 299848 444388 299900 444440
rect 255412 443980 255464 444032
rect 295800 443980 295852 444032
rect 255596 443912 255648 443964
rect 297456 443912 297508 443964
rect 226524 443844 226576 443896
rect 254308 443844 254360 443896
rect 297640 443844 297692 443896
rect 200948 443368 201000 443420
rect 252652 443776 252704 443828
rect 296904 443776 296956 443828
rect 200764 443300 200816 443352
rect 220452 443708 220504 443760
rect 229468 443708 229520 443760
rect 249892 443708 249944 443760
rect 297364 443708 297416 443760
rect 229836 443640 229888 443692
rect 245660 443640 245712 443692
rect 297548 443640 297600 443692
rect 198004 443232 198056 443284
rect 220452 443572 220504 443624
rect 192484 443164 192536 443216
rect 228180 443504 228232 443556
rect 4068 443096 4120 443148
rect 225788 443436 225840 443488
rect 225236 443368 225288 443420
rect 227996 443368 228048 443420
rect 230388 443368 230440 443420
rect 3332 443028 3384 443080
rect 3608 442960 3660 443012
rect 233700 443368 233752 443420
rect 242900 443368 242952 443420
rect 249708 443368 249760 443420
rect 275468 443164 275520 443216
rect 275376 443096 275428 443148
rect 296812 443028 296864 443080
rect 298008 442960 298060 443012
rect 265900 431876 265952 431928
rect 298008 431876 298060 431928
rect 384304 431876 384356 431928
rect 580172 431876 580224 431928
rect 267004 426368 267056 426420
rect 298008 426368 298060 426420
rect 2780 410932 2832 410984
rect 4988 410932 5040 410984
rect 265808 404268 265860 404320
rect 298008 404268 298060 404320
rect 293868 401548 293920 401600
rect 385040 401548 385092 401600
rect 297180 401344 297232 401396
rect 293408 401072 293460 401124
rect 298008 401072 298060 401124
rect 292948 401004 293000 401056
rect 293224 400936 293276 400988
rect 297180 400936 297232 400988
rect 293316 400868 293368 400920
rect 299664 400732 299716 400784
rect 299848 400732 299900 400784
rect 298008 400664 298060 400716
rect 307576 400664 307628 400716
rect 324228 400664 324280 400716
rect 332508 400664 332560 400716
rect 340972 400664 341024 400716
rect 298560 400120 298612 400172
rect 579988 400120 580040 400172
rect 252652 399780 252704 399832
rect 253480 399780 253532 399832
rect 252652 399644 252704 399696
rect 253204 399644 253256 399696
rect 253204 399508 253256 399560
rect 253664 399508 253716 399560
rect 253112 399372 253164 399424
rect 253664 399372 253716 399424
rect 205640 399100 205692 399152
rect 210240 399100 210292 399152
rect 207664 399032 207716 399084
rect 216956 399032 217008 399084
rect 217692 399032 217744 399084
rect 220820 398964 220872 399016
rect 244372 398964 244424 399016
rect 437480 398964 437532 399016
rect 209872 398896 209924 398948
rect 226708 398896 226760 398948
rect 244832 398896 244884 398948
rect 210240 398828 210292 398880
rect 226340 398828 226392 398880
rect 245936 398828 245988 398880
rect 206284 398760 206336 398812
rect 219440 398760 219492 398812
rect 217692 398692 217744 398744
rect 227720 398692 227772 398744
rect 207756 398624 207808 398676
rect 223396 398624 223448 398676
rect 211896 398556 211948 398608
rect 213552 398556 213604 398608
rect 208400 398488 208452 398540
rect 226524 398488 226576 398540
rect 208032 398420 208084 398472
rect 218888 398420 218940 398472
rect 207020 398352 207072 398404
rect 226432 398352 226484 398404
rect 189080 398284 189132 398336
rect 225052 398284 225104 398336
rect 171140 398216 171192 398268
rect 223672 398216 223724 398268
rect 164240 398148 164292 398200
rect 125600 398080 125652 398132
rect 211436 398080 211488 398132
rect 212448 398080 212500 398132
rect 209320 398012 209372 398064
rect 218612 398080 218664 398132
rect 212816 397944 212868 397996
rect 218888 398148 218940 398200
rect 219348 398148 219400 398200
rect 219348 398012 219400 398064
rect 230848 398760 230900 398812
rect 242624 398760 242676 398812
rect 250168 398692 250220 398744
rect 253480 398896 253532 398948
rect 543740 398896 543792 398948
rect 254308 398828 254360 398880
rect 564440 398828 564492 398880
rect 252744 398760 252796 398812
rect 253112 398760 253164 398812
rect 261484 398760 261536 398812
rect 293592 398760 293644 398812
rect 303896 398760 303948 398812
rect 299388 398692 299440 398744
rect 370872 398692 370924 398744
rect 293684 398624 293736 398676
rect 362500 398624 362552 398676
rect 246212 398488 246264 398540
rect 246764 398420 246816 398472
rect 264244 398556 264296 398608
rect 293776 398556 293828 398608
rect 357992 398556 358044 398608
rect 253480 398488 253532 398540
rect 264336 398488 264388 398540
rect 295800 398488 295852 398540
rect 354128 398488 354180 398540
rect 255412 398420 255464 398472
rect 278044 398420 278096 398472
rect 293500 398420 293552 398472
rect 349620 398420 349672 398472
rect 247316 398284 247368 398336
rect 269764 398352 269816 398404
rect 299664 398352 299716 398404
rect 345756 398352 345808 398404
rect 271144 398284 271196 398336
rect 298652 398284 298704 398336
rect 320640 398284 320692 398336
rect 230296 398148 230348 398200
rect 241520 398148 241572 398200
rect 248512 398148 248564 398200
rect 274088 398216 274140 398268
rect 275376 398216 275428 398268
rect 312268 398216 312320 398268
rect 256700 398148 256752 398200
rect 275468 398148 275520 398200
rect 366364 398148 366416 398200
rect 238208 398080 238260 398132
rect 246488 398080 246540 398132
rect 247684 398080 247736 398132
rect 480260 398080 480312 398132
rect 233240 398012 233292 398064
rect 241520 398012 241572 398064
rect 243728 398012 243780 398064
rect 223120 397944 223172 397996
rect 237380 397944 237432 397996
rect 243912 397944 243964 397996
rect 245384 397944 245436 397996
rect 253480 397944 253532 397996
rect 255504 398012 255556 398064
rect 258816 398012 258868 398064
rect 257528 397944 257580 397996
rect 207848 397876 207900 397928
rect 217784 397876 217836 397928
rect 239864 397876 239916 397928
rect 242624 397876 242676 397928
rect 244280 397876 244332 397928
rect 247316 397876 247368 397928
rect 207940 397808 207992 397860
rect 240508 397808 240560 397860
rect 247960 397808 248012 397860
rect 248512 397808 248564 397860
rect 218336 397740 218388 397792
rect 209136 397672 209188 397724
rect 212264 397672 212316 397724
rect 213920 397672 213972 397724
rect 216404 397672 216456 397724
rect 217784 397672 217836 397724
rect 222844 397740 222896 397792
rect 231952 397740 232004 397792
rect 239864 397740 239916 397792
rect 240232 397740 240284 397792
rect 247684 397740 247736 397792
rect 250168 397808 250220 397860
rect 257436 397808 257488 397860
rect 219440 397672 219492 397724
rect 227444 397672 227496 397724
rect 243176 397672 243228 397724
rect 256332 397740 256384 397792
rect 255964 397672 256016 397724
rect 209228 397604 209280 397656
rect 212172 397604 212224 397656
rect 213368 397604 213420 397656
rect 217232 397604 217284 397656
rect 222200 397604 222252 397656
rect 227628 397604 227680 397656
rect 234068 397604 234120 397656
rect 234436 397604 234488 397656
rect 239312 397604 239364 397656
rect 246948 397604 247000 397656
rect 247316 397604 247368 397656
rect 258724 397604 258776 397656
rect 212172 397468 212224 397520
rect 215024 397536 215076 397588
rect 216404 397536 216456 397588
rect 222384 397536 222436 397588
rect 226340 397536 226392 397588
rect 227904 397536 227956 397588
rect 242072 397536 242124 397588
rect 256148 397536 256200 397588
rect 256240 397536 256292 397588
rect 212816 397468 212868 397520
rect 220084 397468 220136 397520
rect 227628 397468 227680 397520
rect 228272 397468 228324 397520
rect 231492 397468 231544 397520
rect 234068 397468 234120 397520
rect 236092 397468 236144 397520
rect 238208 397468 238260 397520
rect 238760 397468 238812 397520
rect 244832 397468 244884 397520
rect 525800 397468 525852 397520
rect 255964 397332 256016 397384
rect 256148 397332 256200 397384
rect 201500 397264 201552 397316
rect 226064 397264 226116 397316
rect 209044 397196 209096 397248
rect 224684 397196 224736 397248
rect 194600 397128 194652 397180
rect 225512 397128 225564 397180
rect 237012 397128 237064 397180
rect 155960 397060 156012 397112
rect 222476 397060 222528 397112
rect 225604 397060 225656 397112
rect 226064 397060 226116 397112
rect 230480 397060 230532 397112
rect 242072 397060 242124 397112
rect 251548 397128 251600 397180
rect 255964 397128 256016 397180
rect 144920 396992 144972 397044
rect 221648 396992 221700 397044
rect 229192 396992 229244 397044
rect 230204 396992 230256 397044
rect 232688 396992 232740 397044
rect 232872 396992 232924 397044
rect 241704 396992 241756 397044
rect 131120 396924 131172 396976
rect 77300 396856 77352 396908
rect 213920 396856 213972 396908
rect 46940 396788 46992 396840
rect 211160 396788 211212 396840
rect 227812 396924 227864 396976
rect 228640 396924 228692 396976
rect 229284 396924 229336 396976
rect 230112 396924 230164 396976
rect 231860 396924 231912 396976
rect 232964 396924 233016 396976
rect 225328 396856 225380 396908
rect 225880 396856 225932 396908
rect 229376 396856 229428 396908
rect 230020 396856 230072 396908
rect 231032 396856 231084 396908
rect 231492 396856 231544 396908
rect 254216 396992 254268 397044
rect 255044 396992 255096 397044
rect 342260 396924 342312 396976
rect 402980 396856 403032 396908
rect 220544 396788 220596 396840
rect 228088 396788 228140 396840
rect 228640 396788 228692 396840
rect 230572 396788 230624 396840
rect 231768 396788 231820 396840
rect 231860 396788 231912 396840
rect 232320 396788 232372 396840
rect 233608 396788 233660 396840
rect 234252 396788 234304 396840
rect 242256 396788 242308 396840
rect 409880 396788 409932 396840
rect 40040 396720 40092 396772
rect 226616 396720 226668 396772
rect 227260 396720 227312 396772
rect 229744 396720 229796 396772
rect 230756 396720 230808 396772
rect 231032 396720 231084 396772
rect 232228 396720 232280 396772
rect 232596 396720 232648 396772
rect 233516 396720 233568 396772
rect 233884 396720 233936 396772
rect 247224 396720 247276 396772
rect 473360 396720 473412 396772
rect 213460 396652 213512 396704
rect 225144 396652 225196 396704
rect 226248 396652 226300 396704
rect 226708 396652 226760 396704
rect 227168 396652 227220 396704
rect 229284 396652 229336 396704
rect 230572 396652 230624 396704
rect 231400 396652 231452 396704
rect 254032 396652 254084 396704
rect 254860 396652 254912 396704
rect 225788 396584 225840 396636
rect 225972 396584 226024 396636
rect 226524 396584 226576 396636
rect 226984 396584 227036 396636
rect 225604 396516 225656 396568
rect 227076 396516 227128 396568
rect 229100 396516 229152 396568
rect 229468 396516 229520 396568
rect 229652 396516 229704 396568
rect 229836 396516 229888 396568
rect 230756 396516 230808 396568
rect 231124 396516 231176 396568
rect 232044 396516 232096 396568
rect 232688 396516 232740 396568
rect 233516 396516 233568 396568
rect 233976 396516 234028 396568
rect 254124 396516 254176 396568
rect 254400 396516 254452 396568
rect 227996 396448 228048 396500
rect 230664 396448 230716 396500
rect 231216 396448 231268 396500
rect 232136 396448 232188 396500
rect 232872 396448 232924 396500
rect 233424 396448 233476 396500
rect 234160 396448 234212 396500
rect 226892 396244 226944 396296
rect 227536 396244 227588 396296
rect 234528 396380 234580 396432
rect 235448 396380 235500 396432
rect 254308 396380 254360 396432
rect 254676 396380 254728 396432
rect 254124 396312 254176 396364
rect 254584 396312 254636 396364
rect 228180 396244 228232 396296
rect 233884 396244 233936 396296
rect 234068 396244 234120 396296
rect 253940 396108 253992 396160
rect 254952 396108 255004 396160
rect 241612 395836 241664 395888
rect 242440 395836 242492 395888
rect 248512 395836 248564 395888
rect 249156 395836 249208 395888
rect 249248 395836 249300 395888
rect 249524 395836 249576 395888
rect 231492 395768 231544 395820
rect 266360 395768 266412 395820
rect 231308 395700 231360 395752
rect 269120 395700 269172 395752
rect 232964 395632 233016 395684
rect 276020 395632 276072 395684
rect 149704 395564 149756 395616
rect 216956 395564 217008 395616
rect 241520 395564 241572 395616
rect 293960 395564 294012 395616
rect 115940 395496 115992 395548
rect 218888 395496 218940 395548
rect 223120 395496 223172 395548
rect 227352 395496 227404 395548
rect 252008 395496 252060 395548
rect 535460 395496 535512 395548
rect 52460 395428 52512 395480
rect 214472 395428 214524 395480
rect 252652 395428 252704 395480
rect 542360 395428 542412 395480
rect 30380 395360 30432 395412
rect 212724 395360 212776 395412
rect 228364 395360 228416 395412
rect 228548 395360 228600 395412
rect 253664 395360 253716 395412
rect 549260 395360 549312 395412
rect 27620 395292 27672 395344
rect 211436 395292 211488 395344
rect 255044 395292 255096 395344
rect 564532 395292 564584 395344
rect 238852 395156 238904 395208
rect 239772 395156 239824 395208
rect 244648 395088 244700 395140
rect 245384 395088 245436 395140
rect 228272 394680 228324 394732
rect 231124 394680 231176 394732
rect 232412 394680 232464 394732
rect 232780 394680 232832 394732
rect 237932 394680 237984 394732
rect 238392 394680 238444 394732
rect 236000 394612 236052 394664
rect 244004 394612 244056 394664
rect 225236 394544 225288 394596
rect 227720 394544 227772 394596
rect 228272 394544 228324 394596
rect 228824 394544 228876 394596
rect 237380 394544 237432 394596
rect 238024 394544 238076 394596
rect 251272 394544 251324 394596
rect 251640 394544 251692 394596
rect 215300 394476 215352 394528
rect 224224 394476 224276 394528
rect 234436 394476 234488 394528
rect 305000 394476 305052 394528
rect 211988 394340 212040 394392
rect 212540 394340 212592 394392
rect 214288 394340 214340 394392
rect 214656 394340 214708 394392
rect 202880 394272 202932 394324
rect 226156 394408 226208 394460
rect 235540 394408 235592 394460
rect 234712 394340 234764 394392
rect 235264 394340 235316 394392
rect 236276 394340 236328 394392
rect 238760 394408 238812 394460
rect 239128 394408 239180 394460
rect 322940 394408 322992 394460
rect 221280 394272 221332 394324
rect 221648 394272 221700 394324
rect 193220 394204 193272 394256
rect 225052 394272 225104 394324
rect 229560 394204 229612 394256
rect 229928 394204 229980 394256
rect 230204 394204 230256 394256
rect 178040 394136 178092 394188
rect 215300 394136 215352 394188
rect 129740 394068 129792 394120
rect 220452 394136 220504 394188
rect 221004 394136 221056 394188
rect 221464 394136 221516 394188
rect 234896 394204 234948 394256
rect 235264 394204 235316 394256
rect 236736 394136 236788 394188
rect 69020 394000 69072 394052
rect 215668 394068 215720 394120
rect 217048 394068 217100 394120
rect 217416 394068 217468 394120
rect 219532 394068 219584 394120
rect 220360 394068 220412 394120
rect 221188 394068 221240 394120
rect 221556 394068 221608 394120
rect 234620 394068 234672 394120
rect 234988 394068 235040 394120
rect 215576 394000 215628 394052
rect 216312 394000 216364 394052
rect 216956 394000 217008 394052
rect 217968 394000 218020 394052
rect 219624 394000 219676 394052
rect 220176 394000 220228 394052
rect 220912 394000 220964 394052
rect 221740 394000 221792 394052
rect 222384 394000 222436 394052
rect 223212 394000 223264 394052
rect 223672 394000 223724 394052
rect 224500 394000 224552 394052
rect 236092 394000 236144 394052
rect 236368 394000 236420 394052
rect 4160 393932 4212 393984
rect 210700 393932 210752 393984
rect 212632 393932 212684 393984
rect 213184 393932 213236 393984
rect 214012 393932 214064 393984
rect 214840 393932 214892 393984
rect 215668 393932 215720 393984
rect 216036 393932 216088 393984
rect 216864 393932 216916 393984
rect 217600 393932 217652 393984
rect 218612 393932 218664 393984
rect 219072 393932 219124 393984
rect 219808 393932 219860 393984
rect 220268 393932 220320 393984
rect 221096 393932 221148 393984
rect 222108 393932 222160 393984
rect 222476 393932 222528 393984
rect 222936 393932 222988 393984
rect 223856 393932 223908 393984
rect 224868 393932 224920 393984
rect 234988 393932 235040 393984
rect 235356 393932 235408 393984
rect 236000 393932 236052 393984
rect 236644 393932 236696 393984
rect 237748 394204 237800 394256
rect 240140 394272 240192 394324
rect 244004 394340 244056 394392
rect 329840 394340 329892 394392
rect 238852 394136 238904 394188
rect 239404 394136 239456 394188
rect 240140 394136 240192 394188
rect 240692 394136 240744 394188
rect 240232 394068 240284 394120
rect 240600 394068 240652 394120
rect 240324 394000 240376 394052
rect 240692 394000 240744 394052
rect 332600 394272 332652 394324
rect 243176 394204 243228 394256
rect 243544 394204 243596 394256
rect 243912 394204 243964 394256
rect 347780 394204 347832 394256
rect 243360 394136 243412 394188
rect 243728 394136 243780 394188
rect 244372 394136 244424 394188
rect 245200 394136 245252 394188
rect 246212 394136 246264 394188
rect 340880 394136 340932 394188
rect 241520 394068 241572 394120
rect 241888 394068 241940 394120
rect 244280 394068 244332 394120
rect 244924 394068 244976 394120
rect 246948 394068 247000 394120
rect 372620 394068 372672 394120
rect 240600 393932 240652 393984
rect 241060 393932 241112 393984
rect 241612 393932 241664 393984
rect 242164 393932 242216 393984
rect 210148 393864 210200 393916
rect 210608 393864 210660 393916
rect 211436 393864 211488 393916
rect 212080 393864 212132 393916
rect 212816 393864 212868 393916
rect 213828 393864 213880 393916
rect 214564 393864 214616 393916
rect 215208 393864 215260 393916
rect 215484 393864 215536 393916
rect 216220 393864 216272 393916
rect 216772 393864 216824 393916
rect 217876 393864 217928 393916
rect 218336 393864 218388 393916
rect 219256 393864 219308 393916
rect 219716 393864 219768 393916
rect 220636 393864 220688 393916
rect 222752 393864 222804 393916
rect 223212 393864 223264 393916
rect 236184 393864 236236 393916
rect 209964 393796 210016 393848
rect 210516 393796 210568 393848
rect 211620 393796 211672 393848
rect 212356 393796 212408 393848
rect 214380 393796 214432 393848
rect 214932 393796 214984 393848
rect 218520 393796 218572 393848
rect 219164 393796 219216 393848
rect 219900 393796 219952 393848
rect 220728 393796 220780 393848
rect 224040 393796 224092 393848
rect 224316 393796 224368 393848
rect 234804 393796 234856 393848
rect 235724 393796 235776 393848
rect 214104 393728 214156 393780
rect 215116 393728 215168 393780
rect 221188 393728 221240 393780
rect 221832 393728 221884 393780
rect 237564 393864 237616 393916
rect 240416 393864 240468 393916
rect 241244 393864 241296 393916
rect 241888 393864 241940 393916
rect 242348 393864 242400 393916
rect 243084 393864 243136 393916
rect 243452 393864 243504 393916
rect 244648 394000 244700 394052
rect 245200 394000 245252 394052
rect 249892 394000 249944 394052
rect 250536 394000 250588 394052
rect 252836 394000 252888 394052
rect 253204 394000 253256 394052
rect 251548 393932 251600 393984
rect 251732 393932 251784 393984
rect 252652 393932 252704 393984
rect 252928 393932 252980 393984
rect 382280 394000 382332 394052
rect 254768 393932 254820 393984
rect 571340 393932 571392 393984
rect 237380 393796 237432 393848
rect 238300 393796 238352 393848
rect 240324 393796 240376 393848
rect 241152 393796 241204 393848
rect 241704 393796 241756 393848
rect 241980 393796 242032 393848
rect 244464 393796 244516 393848
rect 244740 393796 244792 393848
rect 247040 393796 247092 393848
rect 247316 393796 247368 393848
rect 247408 393796 247460 393848
rect 247868 393796 247920 393848
rect 248696 393796 248748 393848
rect 248972 393796 249024 393848
rect 249984 393796 250036 393848
rect 250260 393796 250312 393848
rect 251180 393796 251232 393848
rect 251732 393796 251784 393848
rect 252928 393796 252980 393848
rect 253296 393796 253348 393848
rect 236828 393728 236880 393780
rect 244188 393728 244240 393780
rect 244556 393728 244608 393780
rect 245292 393728 245344 393780
rect 252836 393728 252888 393780
rect 253388 393728 253440 393780
rect 213092 393660 213144 393712
rect 213644 393660 213696 393712
rect 235264 393660 235316 393712
rect 235448 393660 235500 393712
rect 236276 393660 236328 393712
rect 236368 393660 236420 393712
rect 236920 393660 236972 393712
rect 243176 393660 243228 393712
rect 243820 393660 243872 393712
rect 244740 393660 244792 393712
rect 245016 393660 245068 393712
rect 251180 393660 251232 393712
rect 251824 393660 251876 393712
rect 244832 393592 244884 393644
rect 244924 393388 244976 393440
rect 227904 393320 227956 393372
rect 228456 393320 228508 393372
rect 221464 393184 221516 393236
rect 221924 393184 221976 393236
rect 239864 392776 239916 392828
rect 277400 392776 277452 392828
rect 232596 392708 232648 392760
rect 281540 392708 281592 392760
rect 160100 392640 160152 392692
rect 217784 392640 217836 392692
rect 242440 392640 242492 392692
rect 401600 392640 401652 392692
rect 109040 392572 109092 392624
rect 218888 392572 218940 392624
rect 249248 392572 249300 392624
rect 498200 392572 498252 392624
rect 218704 392504 218756 392556
rect 245660 392368 245712 392420
rect 246212 392368 246264 392420
rect 218796 392300 218848 392352
rect 210056 392164 210108 392216
rect 210884 392164 210936 392216
rect 222936 392164 222988 392216
rect 223304 392164 223356 392216
rect 245752 392164 245804 392216
rect 246304 392164 246356 392216
rect 238944 392096 238996 392148
rect 239680 392096 239732 392148
rect 250260 392096 250312 392148
rect 250444 392096 250496 392148
rect 247132 392028 247184 392080
rect 247776 392028 247828 392080
rect 248420 392028 248472 392080
rect 248880 392028 248932 392080
rect 249800 392028 249852 392080
rect 250168 392028 250220 392080
rect 248696 391960 248748 392012
rect 249432 391960 249484 392012
rect 248420 391892 248472 391944
rect 249340 391892 249392 391944
rect 249800 391892 249852 391944
rect 250720 391892 250772 391944
rect 216404 391824 216456 391876
rect 216036 391756 216088 391808
rect 215852 391620 215904 391672
rect 216220 391620 216272 391672
rect 238208 391552 238260 391604
rect 331220 391552 331272 391604
rect 215852 391484 215904 391536
rect 216588 391484 216640 391536
rect 239772 391484 239824 391536
rect 365720 391484 365772 391536
rect 247960 391416 248012 391468
rect 387800 391416 387852 391468
rect 245384 391348 245436 391400
rect 440240 391348 440292 391400
rect 245844 391280 245896 391332
rect 456800 391280 456852 391332
rect 210332 391212 210384 391264
rect 210516 391212 210568 391264
rect 237840 391212 237892 391264
rect 238392 391212 238444 391264
rect 250812 391212 250864 391264
rect 512000 391212 512052 391264
rect 245844 391008 245896 391060
rect 246580 391008 246632 391060
rect 239220 390600 239272 390652
rect 239496 390600 239548 390652
rect 210240 390532 210292 390584
rect 210976 390532 211028 390584
rect 210332 390464 210384 390516
rect 211068 390464 211120 390516
rect 251272 390464 251324 390516
rect 252100 390464 252152 390516
rect 214472 390396 214524 390448
rect 214748 390396 214800 390448
rect 217232 390260 217284 390312
rect 217508 390260 217560 390312
rect 246120 390056 246172 390108
rect 246396 390056 246448 390108
rect 222568 389988 222620 390040
rect 223212 389988 223264 390040
rect 233976 389920 234028 389972
rect 298100 389920 298152 389972
rect 222568 389852 222620 389904
rect 223488 389852 223540 389904
rect 240876 389852 240928 389904
rect 391940 389852 391992 389904
rect 223764 389784 223816 389836
rect 224592 389784 224644 389836
rect 249524 389784 249576 389836
rect 499580 389784 499632 389836
rect 250444 389308 250496 389360
rect 250628 389308 250680 389360
rect 299204 379448 299256 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 98644 372512 98696 372564
rect 295892 365644 295944 365696
rect 580172 365644 580224 365696
rect 106280 363604 106332 363656
rect 209320 363604 209372 363656
rect 2780 358436 2832 358488
rect 4896 358436 4948 358488
rect 92480 355444 92532 355496
rect 217232 355444 217284 355496
rect 232504 355444 232556 355496
rect 284300 355444 284352 355496
rect 42800 355376 42852 355428
rect 213092 355376 213144 355428
rect 244740 355376 244792 355428
rect 445760 355376 445812 355428
rect 37280 355308 37332 355360
rect 213000 355308 213052 355360
rect 250536 355308 250588 355360
rect 514760 355308 514812 355360
rect 169024 354424 169076 354476
rect 218612 354424 218664 354476
rect 88340 354356 88392 354408
rect 213184 354356 213236 354408
rect 91100 354288 91152 354340
rect 217048 354288 217100 354340
rect 231032 354288 231084 354340
rect 262220 354288 262272 354340
rect 86960 354220 87012 354272
rect 217140 354220 217192 354272
rect 246580 354220 246632 354272
rect 357440 354220 357492 354272
rect 70400 354152 70452 354204
rect 212080 354152 212132 354204
rect 240876 354152 240928 354204
rect 393320 354152 393372 354204
rect 60740 354084 60792 354136
rect 211988 354084 212040 354136
rect 228364 354084 228416 354136
rect 232504 354084 232556 354136
rect 245016 354084 245068 354136
rect 440332 354084 440384 354136
rect 62120 354016 62172 354068
rect 214564 354016 214616 354068
rect 229744 354016 229796 354068
rect 240784 354016 240836 354068
rect 251824 354016 251876 354068
rect 534080 354016 534132 354068
rect 56600 353948 56652 354000
rect 214472 353948 214524 354000
rect 229836 353948 229888 354000
rect 244740 353948 244792 354000
rect 253204 353948 253256 354000
rect 546500 353948 546552 354000
rect 299296 353200 299348 353252
rect 580172 353200 580224 353252
rect 198740 352724 198792 352776
rect 225512 352724 225564 352776
rect 180800 352656 180852 352708
rect 224224 352656 224276 352708
rect 235356 352656 235408 352708
rect 316040 352656 316092 352708
rect 160192 352588 160244 352640
rect 223028 352588 223080 352640
rect 240692 352588 240744 352640
rect 385040 352588 385092 352640
rect 5540 352520 5592 352572
rect 210424 352520 210476 352572
rect 243636 352520 243688 352572
rect 423680 352520 423732 352572
rect 225696 351908 225748 351960
rect 226892 351908 226944 351960
rect 238116 351228 238168 351280
rect 357532 351228 357584 351280
rect 85580 351160 85632 351212
rect 210516 351160 210568 351212
rect 254584 351160 254636 351212
rect 572720 351160 572772 351212
rect 110420 340144 110472 340196
rect 208032 340144 208084 340196
rect 23480 338716 23532 338768
rect 209228 338716 209280 338768
rect 258816 334568 258868 334620
rect 581000 334568 581052 334620
rect 24860 333208 24912 333260
rect 209136 333208 209188 333260
rect 258724 333208 258776 333260
rect 436100 333208 436152 333260
rect 296628 325592 296680 325644
rect 580172 325592 580224 325644
rect 3332 320084 3384 320136
rect 199568 320084 199620 320136
rect 296536 313216 296588 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 200948 306280 201000 306332
rect 257528 304240 257580 304292
rect 429200 304240 429252 304292
rect 265716 299412 265768 299464
rect 580172 299412 580224 299464
rect 296444 273164 296496 273216
rect 580172 273164 580224 273216
rect 3148 267656 3200 267708
rect 196716 267656 196768 267708
rect 296352 259360 296404 259412
rect 580172 259360 580224 259412
rect 299112 245556 299164 245608
rect 580172 245556 580224 245608
rect 299020 233180 299072 233232
rect 579988 233180 580040 233232
rect 296260 219376 296312 219428
rect 580172 219376 580224 219428
rect 3056 215228 3108 215280
rect 199476 215228 199528 215280
rect 269856 206932 269908 206984
rect 579804 206932 579856 206984
rect 271236 193128 271288 193180
rect 580172 193128 580224 193180
rect 275284 185580 275336 185632
rect 582380 185580 582432 185632
rect 274088 184152 274140 184204
rect 474740 184152 474792 184204
rect 264336 182792 264388 182844
rect 449900 182792 449952 182844
rect 38660 181432 38712 181484
rect 202144 181432 202196 181484
rect 102232 180072 102284 180124
rect 207940 180072 207992 180124
rect 261484 180072 261536 180124
rect 443000 180072 443052 180124
rect 296168 179324 296220 179376
rect 580172 179324 580224 179376
rect 176660 178712 176712 178764
rect 224132 178712 224184 178764
rect 41420 178644 41472 178696
rect 211896 178644 211948 178696
rect 167000 177556 167052 177608
rect 222936 177556 222988 177608
rect 154580 177488 154632 177540
rect 216036 177488 216088 177540
rect 217048 177488 217100 177540
rect 226708 177488 226760 177540
rect 140780 177420 140832 177472
rect 221556 177420 221608 177472
rect 238024 177420 238076 177472
rect 353300 177420 353352 177472
rect 124220 177352 124272 177404
rect 220084 177352 220136 177404
rect 240600 177352 240652 177404
rect 394700 177352 394752 177404
rect 9680 177284 9732 177336
rect 210332 177284 210384 177336
rect 211528 177284 211580 177336
rect 226800 177284 226852 177336
rect 228272 177284 228324 177336
rect 238024 177284 238076 177336
rect 249064 177284 249116 177336
rect 496820 177284 496872 177336
rect 226892 176672 226944 176724
rect 228180 176672 228232 176724
rect 31760 168988 31812 169040
rect 203708 168988 203760 169040
rect 273996 166948 274048 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 196624 164160 196676 164212
rect 298928 153144 298980 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 192484 150356 192536 150408
rect 295984 139340 296036 139392
rect 580172 139340 580224 139392
rect 268384 126896 268436 126948
rect 580172 126896 580224 126948
rect 298836 113092 298888 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 199384 111732 199436 111784
rect 296076 100648 296128 100700
rect 580172 100648 580224 100700
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 232412 87796 232464 87848
rect 288440 87796 288492 87848
rect 235264 87728 235316 87780
rect 311900 87728 311952 87780
rect 239404 87660 239456 87712
rect 375380 87660 375432 87712
rect 241888 87592 241940 87644
rect 411260 87592 411312 87644
rect 265624 86912 265676 86964
rect 580172 86912 580224 86964
rect 243544 86504 243596 86556
rect 427820 86504 427872 86556
rect 244832 86436 244884 86488
rect 447140 86436 447192 86488
rect 246212 86368 246264 86420
rect 454040 86368 454092 86420
rect 247592 86300 247644 86352
rect 478880 86300 478932 86352
rect 117320 86232 117372 86284
rect 206284 86232 206336 86284
rect 250444 86232 250496 86284
rect 517520 86232 517572 86284
rect 95240 83444 95292 83496
rect 207848 83444 207900 83496
rect 244924 82220 244976 82272
rect 365812 82220 365864 82272
rect 243452 82152 243504 82204
rect 420920 82152 420972 82204
rect 278044 82084 278096 82136
rect 581092 82084 581144 82136
rect 3424 71680 3476 71732
rect 200856 71680 200908 71732
rect 273904 60664 273956 60716
rect 580172 60664 580224 60716
rect 256332 60052 256384 60104
rect 400220 60052 400272 60104
rect 256240 59984 256292 60036
rect 407120 59984 407172 60036
rect 3056 59304 3108 59356
rect 79324 59304 79376 59356
rect 218612 46316 218664 46368
rect 226616 46316 226668 46368
rect 162860 46248 162912 46300
rect 222752 46248 222804 46300
rect 149060 46180 149112 46232
rect 221464 46180 221516 46232
rect 3148 33056 3200 33108
rect 198004 33056 198056 33108
rect 298744 33056 298796 33108
rect 580172 33056 580224 33108
rect 271144 31016 271196 31068
rect 467840 31016 467892 31068
rect 269764 29588 269816 29640
rect 460940 29588 460992 29640
rect 264244 28228 264296 28280
rect 456892 28228 456944 28280
rect 237932 27208 237984 27260
rect 350540 27208 350592 27260
rect 237840 27140 237892 27192
rect 354680 27140 354732 27192
rect 239312 27072 239364 27124
rect 368480 27072 368532 27124
rect 240508 27004 240560 27056
rect 386420 27004 386472 27056
rect 240416 26936 240468 26988
rect 397460 26936 397512 26988
rect 241796 26868 241848 26920
rect 404360 26868 404412 26920
rect 232228 25916 232280 25968
rect 280160 25916 280212 25968
rect 232320 25848 232372 25900
rect 284392 25848 284444 25900
rect 232136 25780 232188 25832
rect 287060 25780 287112 25832
rect 233792 25712 233844 25764
rect 300860 25712 300912 25764
rect 235172 25644 235224 25696
rect 318800 25644 318852 25696
rect 236460 25576 236512 25628
rect 336740 25576 336792 25628
rect 255412 25508 255464 25560
rect 578240 25508 578292 25560
rect 250352 24420 250404 24472
rect 510620 24420 510672 24472
rect 250260 24352 250312 24404
rect 514852 24352 514904 24404
rect 251732 24284 251784 24336
rect 524420 24284 524472 24336
rect 251640 24216 251692 24268
rect 528560 24216 528612 24268
rect 251548 24148 251600 24200
rect 531320 24148 531372 24200
rect 254492 24080 254544 24132
rect 567200 24080 567252 24132
rect 246028 23128 246080 23180
rect 459560 23128 459612 23180
rect 246120 23060 246172 23112
rect 463700 23060 463752 23112
rect 247500 22992 247552 23044
rect 477500 22992 477552 23044
rect 247408 22924 247460 22976
rect 481640 22924 481692 22976
rect 248880 22856 248932 22908
rect 490012 22856 490064 22908
rect 248972 22788 249024 22840
rect 492680 22788 492732 22840
rect 250168 22720 250220 22772
rect 506572 22720 506624 22772
rect 240324 21632 240376 21684
rect 396080 21632 396132 21684
rect 241704 21564 241756 21616
rect 407212 21564 407264 21616
rect 244648 21496 244700 21548
rect 438860 21496 438912 21548
rect 244464 21428 244516 21480
rect 441620 21428 441672 21480
rect 244556 21360 244608 21412
rect 448520 21360 448572 21412
rect 3424 20612 3476 20664
rect 200764 20612 200816 20664
rect 235080 20272 235132 20324
rect 317420 20272 317472 20324
rect 234988 20204 235040 20256
rect 321560 20204 321612 20256
rect 237748 20136 237800 20188
rect 349160 20136 349212 20188
rect 239128 20068 239180 20120
rect 367100 20068 367152 20120
rect 239036 20000 239088 20052
rect 371240 20000 371292 20052
rect 239220 19932 239272 19984
rect 374000 19932 374052 19984
rect 232044 18912 232096 18964
rect 285680 18912 285732 18964
rect 233608 18844 233660 18896
rect 296720 18844 296772 18896
rect 233700 18776 233752 18828
rect 299572 18776 299624 18828
rect 233516 18708 233568 18760
rect 303620 18708 303672 18760
rect 234896 18640 234948 18692
rect 314660 18640 314712 18692
rect 247316 18572 247368 18624
rect 471980 18572 472032 18624
rect 233884 17620 233936 17672
rect 271880 17620 271932 17672
rect 231952 17552 232004 17604
rect 278780 17552 278832 17604
rect 231860 17484 231912 17536
rect 282920 17484 282972 17536
rect 240232 17416 240284 17468
rect 389180 17416 389232 17468
rect 254400 17348 254452 17400
rect 563060 17348 563112 17400
rect 254216 17280 254268 17332
rect 565820 17280 565872 17332
rect 254308 17212 254360 17264
rect 569960 17212 570012 17264
rect 251456 16124 251508 16176
rect 527824 16124 527876 16176
rect 251364 16056 251416 16108
rect 531412 16056 531464 16108
rect 253112 15988 253164 16040
rect 545488 15988 545540 16040
rect 114008 15920 114060 15972
rect 218520 15920 218572 15972
rect 253020 15920 253072 15972
rect 548616 15920 548668 15972
rect 35992 15852 36044 15904
rect 212908 15852 212960 15904
rect 252928 15852 252980 15904
rect 552664 15852 552716 15904
rect 123024 14900 123076 14952
rect 219992 14900 220044 14952
rect 256148 14900 256200 14952
rect 422576 14900 422628 14952
rect 105728 14832 105780 14884
rect 218428 14832 218480 14884
rect 248604 14832 248656 14884
rect 492312 14832 492364 14884
rect 98184 14764 98236 14816
rect 216956 14764 217008 14816
rect 248788 14764 248840 14816
rect 495440 14764 495492 14816
rect 75000 14696 75052 14748
rect 215944 14696 215996 14748
rect 248512 14696 248564 14748
rect 498936 14696 498988 14748
rect 44180 14628 44232 14680
rect 212816 14628 212868 14680
rect 248696 14628 248748 14680
rect 502984 14628 503036 14680
rect 34520 14560 34572 14612
rect 211804 14560 211856 14612
rect 250076 14560 250128 14612
rect 509608 14560 509660 14612
rect 22560 14492 22612 14544
rect 211436 14492 211488 14544
rect 249984 14492 250036 14544
rect 513380 14492 513432 14544
rect 17960 14424 18012 14476
rect 211344 14424 211396 14476
rect 249892 14424 249944 14476
rect 517152 14424 517204 14476
rect 80888 13540 80940 13592
rect 215852 13540 215904 13592
rect 77392 13472 77444 13524
rect 215576 13472 215628 13524
rect 243360 13472 243412 13524
rect 425704 13472 425756 13524
rect 73344 13404 73396 13456
rect 215668 13404 215720 13456
rect 245936 13404 245988 13456
rect 459192 13404 459244 13456
rect 69848 13336 69900 13388
rect 215760 13336 215812 13388
rect 245752 13336 245804 13388
rect 462320 13336 462372 13388
rect 59360 13268 59412 13320
rect 214380 13268 214432 13320
rect 245844 13268 245896 13320
rect 465816 13268 465868 13320
rect 56048 13200 56100 13252
rect 214288 13200 214340 13252
rect 247040 13200 247092 13252
rect 473452 13200 473504 13252
rect 8760 13132 8812 13184
rect 210240 13132 210292 13184
rect 247224 13132 247276 13184
rect 476488 13132 476540 13184
rect 3608 13064 3660 13116
rect 210148 13064 210200 13116
rect 247132 13064 247184 13116
rect 481732 13064 481784 13116
rect 240140 12112 240192 12164
rect 390652 12112 390704 12164
rect 15936 12044 15988 12096
rect 178684 12044 178736 12096
rect 178776 12044 178828 12096
rect 214196 12044 214248 12096
rect 243268 12044 243320 12096
rect 423772 12044 423824 12096
rect 44272 11976 44324 12028
rect 213276 11976 213328 12028
rect 243084 11976 243136 12028
rect 426808 11976 426860 12028
rect 36728 11908 36780 11960
rect 212632 11908 212684 11960
rect 243176 11908 243228 11960
rect 430856 11908 430908 11960
rect 33600 11840 33652 11892
rect 212724 11840 212776 11892
rect 244280 11840 244332 11892
rect 445024 11840 445076 11892
rect 26240 11772 26292 11824
rect 211620 11772 211672 11824
rect 244372 11772 244424 11824
rect 448612 11772 448664 11824
rect 21824 11704 21876 11756
rect 212356 11704 212408 11756
rect 245660 11704 245712 11756
rect 455696 11704 455748 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 171784 10752 171836 10804
rect 218336 10752 218388 10804
rect 111616 10684 111668 10736
rect 218704 10684 218756 10736
rect 108120 10616 108172 10668
rect 218796 10616 218848 10668
rect 238852 10616 238904 10668
rect 374092 10616 374144 10668
rect 104072 10548 104124 10600
rect 218244 10548 218296 10600
rect 247684 10548 247736 10600
rect 384304 10548 384356 10600
rect 97448 10480 97500 10532
rect 216772 10480 216824 10532
rect 242440 10480 242492 10532
rect 379520 10480 379572 10532
rect 93952 10412 94004 10464
rect 216864 10412 216916 10464
rect 238944 10412 238996 10464
rect 377680 10412 377732 10464
rect 89904 10344 89956 10396
rect 217416 10344 217468 10396
rect 241520 10344 241572 10396
rect 406016 10344 406068 10396
rect 11152 10276 11204 10328
rect 188344 10276 188396 10328
rect 241612 10276 241664 10328
rect 409144 10276 409196 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 79692 9324 79744 9376
rect 216128 9324 216180 9376
rect 76196 9256 76248 9308
rect 215484 9256 215536 9308
rect 237656 9256 237708 9308
rect 349252 9256 349304 9308
rect 72608 9188 72660 9240
rect 216220 9188 216272 9240
rect 237564 9188 237616 9240
rect 352840 9188 352892 9240
rect 62028 9120 62080 9172
rect 214104 9120 214156 9172
rect 237472 9120 237524 9172
rect 356336 9120 356388 9172
rect 58440 9052 58492 9104
rect 214012 9052 214064 9104
rect 237380 9052 237432 9104
rect 359924 9052 359976 9104
rect 7656 8984 7708 9036
rect 210056 8984 210108 9036
rect 238760 8984 238812 9036
rect 370596 8984 370648 9036
rect 2872 8916 2924 8968
rect 209964 8916 210016 8968
rect 257436 8916 257488 8968
rect 415492 8916 415544 8968
rect 197912 7964 197964 8016
rect 225420 7964 225472 8016
rect 158904 7896 158956 7948
rect 222660 7896 222712 7948
rect 151912 7828 151964 7880
rect 221096 7828 221148 7880
rect 148324 7760 148376 7812
rect 221188 7760 221240 7812
rect 233424 7760 233476 7812
rect 306748 7760 306800 7812
rect 144736 7692 144788 7744
rect 221280 7692 221332 7744
rect 234712 7692 234764 7744
rect 320916 7692 320968 7744
rect 142436 7624 142488 7676
rect 221372 7624 221424 7676
rect 234804 7624 234856 7676
rect 324412 7624 324464 7676
rect 54944 7556 54996 7608
rect 214748 7556 214800 7608
rect 252836 7556 252888 7608
rect 553768 7556 553820 7608
rect 230756 6808 230808 6860
rect 267740 6808 267792 6860
rect 230664 6740 230716 6792
rect 268844 6740 268896 6792
rect 234620 6672 234672 6724
rect 317328 6672 317380 6724
rect 200304 6604 200356 6656
rect 225328 6604 225380 6656
rect 236276 6604 236328 6656
rect 332692 6604 332744 6656
rect 187332 6536 187384 6588
rect 223856 6536 223908 6588
rect 236184 6536 236236 6588
rect 336280 6536 336332 6588
rect 183744 6468 183796 6520
rect 223764 6468 223816 6520
rect 236368 6468 236420 6520
rect 342168 6468 342220 6520
rect 180248 6400 180300 6452
rect 224040 6400 224092 6452
rect 242900 6400 242952 6452
rect 418988 6400 419040 6452
rect 176752 6332 176804 6384
rect 223948 6332 224000 6384
rect 242992 6332 243044 6384
rect 420184 6332 420236 6384
rect 169576 6264 169628 6316
rect 222568 6264 222620 6316
rect 256056 6264 256108 6316
rect 562048 6264 562100 6316
rect 134156 6196 134208 6248
rect 219900 6196 219952 6248
rect 254124 6196 254176 6248
rect 569132 6196 569184 6248
rect 128176 6128 128228 6180
rect 219808 6128 219860 6180
rect 254032 6128 254084 6180
rect 572720 6128 572772 6180
rect 230940 6060 230992 6112
rect 265348 6060 265400 6112
rect 230848 5992 230900 6044
rect 261760 5992 261812 6044
rect 201592 5380 201644 5432
rect 225788 5380 225840 5432
rect 196808 5312 196860 5364
rect 225880 5312 225932 5364
rect 166080 5244 166132 5296
rect 222384 5244 222436 5296
rect 150624 5176 150676 5228
rect 147128 5108 147180 5160
rect 162492 5176 162544 5228
rect 222476 5176 222528 5228
rect 249800 5176 249852 5228
rect 519544 5176 519596 5228
rect 157800 5108 157852 5160
rect 223212 5108 223264 5160
rect 251180 5108 251232 5160
rect 533712 5108 533764 5160
rect 221648 5040 221700 5092
rect 251272 5040 251324 5092
rect 537208 5040 537260 5092
rect 220912 4972 220964 5024
rect 252652 4972 252704 5024
rect 547880 4972 547932 5024
rect 143540 4904 143592 4956
rect 221004 4904 221056 4956
rect 229468 4904 229520 4956
rect 241704 4904 241756 4956
rect 252560 4904 252612 4956
rect 551468 4904 551520 4956
rect 132960 4836 133012 4888
rect 219716 4836 219768 4888
rect 229652 4836 229704 4888
rect 251180 4836 251232 4888
rect 252744 4836 252796 4888
rect 554964 4836 555016 4888
rect 19432 4768 19484 4820
rect 203524 4768 203576 4820
rect 205088 4768 205140 4820
rect 225144 4768 225196 4820
rect 229560 4768 229612 4820
rect 252376 4768 252428 4820
rect 254952 4768 255004 4820
rect 560852 4768 560904 4820
rect 228088 4088 228140 4140
rect 229836 4088 229888 4140
rect 230572 4088 230624 4140
rect 239404 4088 239456 4140
rect 242164 4088 242216 4140
rect 259460 4088 259512 4140
rect 217968 4020 218020 4072
rect 223948 4020 224000 4072
rect 231768 4020 231820 4072
rect 95148 3952 95200 4004
rect 149704 3952 149756 4004
rect 219256 3952 219308 4004
rect 222844 3952 222896 4004
rect 227904 3952 227956 4004
rect 233424 3952 233476 4004
rect 234896 4020 234948 4072
rect 258264 4020 258316 4072
rect 260656 3952 260708 4004
rect 115204 3884 115256 3936
rect 171784 3884 171836 3936
rect 186136 3884 186188 3936
rect 224316 3884 224368 3936
rect 227996 3884 228048 3936
rect 235816 3884 235868 3936
rect 236092 3884 236144 3936
rect 239312 3884 239364 3936
rect 239404 3884 239456 3936
rect 271236 3884 271288 3936
rect 112812 3816 112864 3868
rect 169024 3816 169076 3868
rect 184940 3816 184992 3868
rect 209044 3816 209096 3868
rect 219348 3816 219400 3868
rect 264152 3816 264204 3868
rect 284300 3816 284352 3868
rect 285036 3816 285088 3868
rect 82084 3748 82136 3800
rect 138664 3748 138716 3800
rect 151820 3748 151872 3800
rect 153016 3748 153068 3800
rect 168380 3748 168432 3800
rect 207756 3748 207808 3800
rect 215668 3748 215720 3800
rect 225604 3748 225656 3800
rect 233332 3748 233384 3800
rect 296076 3748 296128 3800
rect 118792 3680 118844 3732
rect 185584 3680 185636 3732
rect 214472 3680 214524 3732
rect 226524 3680 226576 3732
rect 234252 3680 234304 3732
rect 299664 3680 299716 3732
rect 135352 3612 135404 3664
rect 207664 3612 207716 3664
rect 213368 3612 213420 3664
rect 227444 3612 227496 3664
rect 229008 3612 229060 3664
rect 237012 3612 237064 3664
rect 239496 3612 239548 3664
rect 335084 3612 335136 3664
rect 12348 3544 12400 3596
rect 88248 3544 88300 3596
rect 88984 3544 89036 3596
rect 129372 3544 129424 3596
rect 219532 3544 219584 3596
rect 229376 3544 229428 3596
rect 13544 3476 13596 3528
rect 118700 3476 118752 3528
rect 119896 3476 119948 3528
rect 126980 3476 127032 3528
rect 219624 3476 219676 3528
rect 231124 3476 231176 3528
rect 232228 3476 232280 3528
rect 236552 3476 236604 3528
rect 44180 3408 44232 3460
rect 45100 3408 45152 3460
rect 52552 3408 52604 3460
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 135260 3340 135312 3392
rect 136456 3340 136508 3392
rect 176660 3408 176712 3460
rect 177856 3408 177908 3460
rect 182548 3408 182600 3460
rect 223672 3408 223724 3460
rect 229192 3408 229244 3460
rect 246396 3544 246448 3596
rect 257344 3544 257396 3596
rect 465172 3544 465224 3596
rect 473360 3544 473412 3596
rect 474188 3544 474240 3596
rect 481640 3544 481692 3596
rect 482468 3544 482520 3596
rect 489920 3544 489972 3596
rect 490748 3544 490800 3596
rect 239404 3476 239456 3528
rect 247592 3476 247644 3528
rect 248420 3476 248472 3528
rect 501788 3476 501840 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 581000 3476 581052 3528
rect 581828 3476 581880 3528
rect 255964 3408 256016 3460
rect 530124 3408 530176 3460
rect 178776 3340 178828 3392
rect 201500 3340 201552 3392
rect 202696 3340 202748 3392
rect 221556 3340 221608 3392
rect 225696 3340 225748 3392
rect 230112 3340 230164 3392
rect 244096 3340 244148 3392
rect 299572 3340 299624 3392
rect 300768 3340 300820 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 456892 3340 456944 3392
rect 458088 3340 458140 3392
rect 229284 3272 229336 3324
rect 20628 3204 20680 3256
rect 25504 3204 25556 3256
rect 236552 3272 236604 3324
rect 239404 3272 239456 3324
rect 240784 3272 240836 3324
rect 232504 3068 232556 3120
rect 234620 3068 234672 3120
rect 248788 3204 248840 3256
rect 236644 3136 236696 3188
rect 242900 3136 242952 3188
rect 249984 3068 250036 3120
rect 227628 2864 227680 2916
rect 231032 2864 231084 2916
rect 423680 1368 423732 1420
rect 424968 1368 425020 1420
rect 448520 1368 448572 1420
rect 449808 1368 449860 1420
rect 365720 1096 365772 1148
rect 367008 1096 367060 1148
rect 390560 1096 390612 1148
rect 391848 1096 391900 1148
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3344 565894 3372 566879
rect 3332 565888 3384 565894
rect 3332 565830 3384 565836
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553450 3188 553823
rect 3148 553444 3200 553450
rect 3148 553386 3200 553392
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3252 474774 3280 475623
rect 3240 474768 3292 474774
rect 3240 474710 3292 474716
rect 2870 462632 2926 462641
rect 2870 462567 2926 462576
rect 2884 462398 2912 462567
rect 2872 462392 2924 462398
rect 2872 462334 2924 462340
rect 3238 449576 3294 449585
rect 3238 449511 3294 449520
rect 3252 447846 3280 449511
rect 3436 448050 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 449886 3556 671191
rect 3606 658200 3662 658209
rect 3606 658135 3662 658144
rect 3516 449880 3568 449886
rect 3516 449822 3568 449828
rect 3424 448044 3476 448050
rect 3424 447986 3476 447992
rect 3620 447982 3648 658135
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3712 448186 3740 632023
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3700 448180 3752 448186
rect 3700 448122 3752 448128
rect 3608 447976 3660 447982
rect 3608 447918 3660 447924
rect 3804 447914 3832 619103
rect 3882 606112 3938 606121
rect 3882 606047 3938 606056
rect 3896 449206 3924 606047
rect 3974 580000 4030 580009
rect 3974 579935 4030 579944
rect 3884 449200 3936 449206
rect 3884 449142 3936 449148
rect 3988 448118 4016 579935
rect 4066 514856 4122 514865
rect 4066 514791 4122 514800
rect 4080 464438 4108 514791
rect 4068 464432 4120 464438
rect 4068 464374 4120 464380
rect 6932 457502 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 22744 553444 22796 553450
rect 22744 553386 22796 553392
rect 14464 527196 14516 527202
rect 14464 527138 14516 527144
rect 10324 501016 10376 501022
rect 10324 500958 10376 500964
rect 10336 469946 10364 500958
rect 10324 469940 10376 469946
rect 10324 469882 10376 469888
rect 14476 460290 14504 527138
rect 22756 468518 22784 553386
rect 22744 468512 22796 468518
rect 22744 468454 22796 468460
rect 14464 460284 14516 460290
rect 14464 460226 14516 460232
rect 6920 457496 6972 457502
rect 6920 457438 6972 457444
rect 23492 448526 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 32404 565888 32456 565894
rect 32404 565830 32456 565836
rect 32416 472734 32444 565830
rect 32404 472728 32456 472734
rect 32404 472670 32456 472676
rect 40052 458862 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40684 474768 40736 474774
rect 40684 474710 40736 474716
rect 40696 471306 40724 474710
rect 40684 471300 40736 471306
rect 40684 471242 40736 471248
rect 71792 461718 71820 702986
rect 89180 700330 89208 703520
rect 105464 700398 105492 703520
rect 137848 700466 137876 703520
rect 154132 700534 154160 703520
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 170324 699718 170352 703520
rect 182824 700528 182876 700534
rect 182824 700470 182876 700476
rect 178684 700460 178736 700466
rect 178684 700402 178736 700408
rect 174544 700392 174596 700398
rect 174544 700334 174596 700340
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171784 699712 171836 699718
rect 171784 699654 171836 699660
rect 78586 636440 78642 636449
rect 78586 636375 78642 636384
rect 78310 635352 78366 635361
rect 78310 635287 78366 635296
rect 78218 633720 78274 633729
rect 78218 633655 78274 633664
rect 77758 632632 77814 632641
rect 77758 632567 77814 632576
rect 77772 523569 77800 632567
rect 78126 631000 78182 631009
rect 78126 630935 78182 630944
rect 77850 629640 77906 629649
rect 77850 629575 77906 629584
rect 77758 523560 77814 523569
rect 77758 523495 77814 523504
rect 77666 520976 77722 520985
rect 77666 520911 77722 520920
rect 77680 489802 77708 520911
rect 77668 489796 77720 489802
rect 77668 489738 77720 489744
rect 77772 489530 77800 523495
rect 77864 521665 77892 629575
rect 78034 628008 78090 628017
rect 78034 627943 78090 627952
rect 77942 608696 77998 608705
rect 77942 608631 77998 608640
rect 77850 521656 77906 521665
rect 77850 521591 77906 521600
rect 77956 498681 77984 608631
rect 78048 599962 78076 627943
rect 78140 600030 78168 630935
rect 78128 600024 78180 600030
rect 78128 599966 78180 599972
rect 78036 599956 78088 599962
rect 78036 599898 78088 599904
rect 78232 599826 78260 633655
rect 78220 599820 78272 599826
rect 78220 599762 78272 599768
rect 78324 584458 78352 635287
rect 78402 610056 78458 610065
rect 78402 609991 78458 610000
rect 78416 599690 78444 609991
rect 78494 607744 78550 607753
rect 78494 607679 78550 607688
rect 78508 599758 78536 607679
rect 78600 599894 78628 636375
rect 78588 599888 78640 599894
rect 78588 599830 78640 599836
rect 78496 599752 78548 599758
rect 78496 599694 78548 599700
rect 78404 599684 78456 599690
rect 78404 599626 78456 599632
rect 102874 597544 102930 597553
rect 102874 597479 102930 597488
rect 111706 597544 111762 597553
rect 111706 597479 111762 597488
rect 92478 597408 92534 597417
rect 92478 597343 92534 597352
rect 100666 597408 100722 597417
rect 100666 597343 100722 597352
rect 92492 596358 92520 597343
rect 99286 597272 99342 597281
rect 99286 597207 99342 597216
rect 94042 597136 94098 597145
rect 99300 597106 99328 597207
rect 100680 597174 100708 597343
rect 102888 597310 102916 597479
rect 102876 597304 102928 597310
rect 102876 597246 102928 597252
rect 104806 597272 104862 597281
rect 104806 597207 104808 597216
rect 104860 597207 104862 597216
rect 104808 597178 104860 597184
rect 100668 597168 100720 597174
rect 100668 597110 100720 597116
rect 102046 597136 102102 597145
rect 94042 597071 94098 597080
rect 99288 597100 99340 597106
rect 79784 596352 79836 596358
rect 79784 596294 79836 596300
rect 92480 596352 92532 596358
rect 92480 596294 92532 596300
rect 78312 584452 78364 584458
rect 78312 584394 78364 584400
rect 78324 526561 78352 584394
rect 78494 526688 78550 526697
rect 78494 526623 78550 526632
rect 78310 526552 78366 526561
rect 78310 526487 78366 526496
rect 78310 523696 78366 523705
rect 78310 523631 78366 523640
rect 78126 521656 78182 521665
rect 78126 521591 78182 521600
rect 78140 520305 78168 521591
rect 78126 520296 78182 520305
rect 78126 520231 78182 520240
rect 78034 499896 78090 499905
rect 78034 499831 78090 499840
rect 77942 498672 77998 498681
rect 77942 498607 77998 498616
rect 77760 489524 77812 489530
rect 77760 489466 77812 489472
rect 77956 475454 77984 498607
rect 78048 489462 78076 499831
rect 78140 489598 78168 520231
rect 78324 489666 78352 523631
rect 78402 498400 78458 498409
rect 78402 498335 78458 498344
rect 78416 489734 78444 498335
rect 78508 489870 78536 526623
rect 78586 517984 78642 517993
rect 78586 517919 78642 517928
rect 78496 489864 78548 489870
rect 78496 489806 78548 489812
rect 78404 489728 78456 489734
rect 78404 489670 78456 489676
rect 78312 489660 78364 489666
rect 78312 489602 78364 489608
rect 78128 489592 78180 489598
rect 78128 489534 78180 489540
rect 78036 489456 78088 489462
rect 78036 489398 78088 489404
rect 78600 489394 78628 517919
rect 78588 489388 78640 489394
rect 78588 489330 78640 489336
rect 79796 488510 79824 596294
rect 94056 596290 94084 597071
rect 102046 597071 102102 597080
rect 99288 597042 99340 597048
rect 102060 597038 102088 597071
rect 102048 597032 102100 597038
rect 102048 596974 102100 596980
rect 103426 597000 103482 597009
rect 103426 596935 103482 596944
rect 106186 597000 106242 597009
rect 106186 596935 106188 596944
rect 103440 596902 103468 596935
rect 106240 596935 106242 596944
rect 106188 596906 106240 596912
rect 103428 596896 103480 596902
rect 97906 596864 97962 596873
rect 103428 596838 103480 596844
rect 97906 596799 97908 596808
rect 97960 596799 97962 596808
rect 97908 596770 97960 596776
rect 95238 596320 95294 596329
rect 79968 596284 80020 596290
rect 79968 596226 80020 596232
rect 94044 596284 94096 596290
rect 95238 596255 95294 596264
rect 94044 596226 94096 596232
rect 79876 596216 79928 596222
rect 79876 596158 79928 596164
rect 79784 488504 79836 488510
rect 79784 488446 79836 488452
rect 79888 488374 79916 596158
rect 79980 488442 80008 596226
rect 95252 596222 95280 596255
rect 95240 596216 95292 596222
rect 95240 596158 95292 596164
rect 111720 581670 111748 597479
rect 131026 597000 131082 597009
rect 131026 596935 131082 596944
rect 126886 596728 126942 596737
rect 126886 596663 126942 596672
rect 126900 596358 126928 596663
rect 131040 596426 131068 596935
rect 136546 596592 136602 596601
rect 136546 596527 136602 596536
rect 140686 596592 140742 596601
rect 140686 596527 140688 596536
rect 136560 596494 136588 596527
rect 140740 596527 140742 596536
rect 140688 596498 140740 596504
rect 136548 596488 136600 596494
rect 136548 596430 136600 596436
rect 131028 596420 131080 596426
rect 131028 596362 131080 596368
rect 126888 596352 126940 596358
rect 115846 596320 115902 596329
rect 115846 596255 115902 596264
rect 121366 596320 121422 596329
rect 126888 596294 126940 596300
rect 121366 596255 121368 596264
rect 115860 596222 115888 596255
rect 121420 596255 121422 596264
rect 121368 596226 121420 596232
rect 115848 596216 115900 596222
rect 115848 596158 115900 596164
rect 111708 581664 111760 581670
rect 111708 581606 111760 581612
rect 92940 488504 92992 488510
rect 92938 488472 92940 488481
rect 92992 488472 92994 488481
rect 79968 488436 80020 488442
rect 92938 488407 92994 488416
rect 94226 488472 94282 488481
rect 94226 488407 94228 488416
rect 79968 488378 80020 488384
rect 94280 488407 94282 488416
rect 95330 488472 95386 488481
rect 95330 488407 95386 488416
rect 97814 488472 97870 488481
rect 97814 488407 97870 488416
rect 98918 488472 98974 488481
rect 98918 488407 98974 488416
rect 100022 488472 100078 488481
rect 100022 488407 100078 488416
rect 101126 488472 101182 488481
rect 101126 488407 101182 488416
rect 102414 488472 102470 488481
rect 102414 488407 102470 488416
rect 104806 488472 104862 488481
rect 104806 488407 104862 488416
rect 105726 488472 105782 488481
rect 105726 488407 105782 488416
rect 94228 488378 94280 488384
rect 95344 488374 95372 488407
rect 79876 488368 79928 488374
rect 79876 488310 79928 488316
rect 95332 488368 95384 488374
rect 95332 488310 95384 488316
rect 97828 487490 97856 488407
rect 97816 487484 97868 487490
rect 97816 487426 97868 487432
rect 98932 487354 98960 488407
rect 98920 487348 98972 487354
rect 98920 487290 98972 487296
rect 100036 487218 100064 488407
rect 101140 487830 101168 488407
rect 101128 487824 101180 487830
rect 101128 487766 101180 487772
rect 102428 487422 102456 488407
rect 104820 487966 104848 488407
rect 105740 488034 105768 488407
rect 105818 488200 105874 488209
rect 105818 488135 105874 488144
rect 111706 488200 111762 488209
rect 111706 488135 111762 488144
rect 105728 488028 105780 488034
rect 105728 487970 105780 487976
rect 104808 487960 104860 487966
rect 103426 487928 103482 487937
rect 104808 487902 104860 487908
rect 103426 487863 103428 487872
rect 103480 487863 103482 487872
rect 103428 487834 103480 487840
rect 102416 487416 102468 487422
rect 102416 487358 102468 487364
rect 100024 487212 100076 487218
rect 100024 487154 100076 487160
rect 105832 482390 105860 488135
rect 105820 482384 105872 482390
rect 105820 482326 105872 482332
rect 77944 475448 77996 475454
rect 77944 475390 77996 475396
rect 71780 461712 71832 461718
rect 71780 461654 71832 461660
rect 40040 458856 40092 458862
rect 40040 458798 40092 458804
rect 111720 449274 111748 488135
rect 115846 487248 115902 487257
rect 115846 487183 115902 487192
rect 121366 487248 121422 487257
rect 121366 487183 121422 487192
rect 126886 487248 126942 487257
rect 126886 487183 126942 487192
rect 131026 487248 131082 487257
rect 131026 487183 131082 487192
rect 136546 487248 136602 487257
rect 136546 487183 136602 487192
rect 140686 487248 140742 487257
rect 140686 487183 140742 487192
rect 115860 449342 115888 487183
rect 121380 467158 121408 487183
rect 126900 479738 126928 487183
rect 126888 479732 126940 479738
rect 126888 479674 126940 479680
rect 121368 467152 121420 467158
rect 121368 467094 121420 467100
rect 131040 461786 131068 487183
rect 136560 465866 136588 487183
rect 136548 465860 136600 465866
rect 136548 465802 136600 465808
rect 131028 461780 131080 461786
rect 131028 461722 131080 461728
rect 140700 449410 140728 487183
rect 171796 451994 171824 699654
rect 173162 596864 173218 596873
rect 173162 596799 173218 596808
rect 172152 596556 172204 596562
rect 172152 596498 172204 596504
rect 171876 596420 171928 596426
rect 171876 596362 171928 596368
rect 171784 451988 171836 451994
rect 171784 451930 171836 451936
rect 140688 449404 140740 449410
rect 140688 449346 140740 449352
rect 115848 449336 115900 449342
rect 115848 449278 115900 449284
rect 111708 449268 111760 449274
rect 111708 449210 111760 449216
rect 171888 449002 171916 596362
rect 171968 596284 172020 596290
rect 171968 596226 172020 596232
rect 171980 458930 172008 596226
rect 172060 596216 172112 596222
rect 172060 596158 172112 596164
rect 172072 478310 172100 596158
rect 172164 485178 172192 596498
rect 172152 485172 172204 485178
rect 172152 485114 172204 485120
rect 172060 478304 172112 478310
rect 172060 478246 172112 478252
rect 173176 474162 173204 596799
rect 173348 596488 173400 596494
rect 173348 596430 173400 596436
rect 173256 596352 173308 596358
rect 173256 596294 173308 596300
rect 173268 481166 173296 596294
rect 173360 489258 173388 596430
rect 173348 489252 173400 489258
rect 173348 489194 173400 489200
rect 173256 481160 173308 481166
rect 173256 481102 173308 481108
rect 173164 474156 173216 474162
rect 173164 474098 173216 474104
rect 171968 458924 172020 458930
rect 171968 458866 172020 458872
rect 174556 457570 174584 700334
rect 178696 467294 178724 700402
rect 178684 467288 178736 467294
rect 178684 467230 178736 467236
rect 174544 457564 174596 457570
rect 174544 457506 174596 457512
rect 182836 453490 182864 700470
rect 202800 700466 202828 703520
rect 188896 700460 188948 700466
rect 188896 700402 188948 700408
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 184204 700324 184256 700330
rect 184204 700266 184256 700272
rect 188804 700324 188856 700330
rect 188804 700266 188856 700272
rect 182824 453484 182876 453490
rect 182824 453426 182876 453432
rect 171876 448996 171928 449002
rect 171876 448938 171928 448944
rect 23480 448520 23532 448526
rect 23480 448462 23532 448468
rect 184216 448254 184244 700266
rect 187330 637120 187386 637129
rect 187330 637055 187386 637064
rect 186778 636032 186834 636041
rect 186778 635967 186834 635976
rect 186792 584458 186820 635967
rect 186870 634400 186926 634409
rect 186870 634335 186926 634344
rect 186884 599826 186912 634335
rect 187238 631680 187294 631689
rect 187238 631615 187294 631624
rect 187146 628688 187202 628697
rect 187146 628623 187202 628632
rect 187054 610328 187110 610337
rect 187054 610263 187110 610272
rect 186962 608424 187018 608433
rect 186962 608359 187018 608368
rect 186872 599820 186924 599826
rect 186872 599762 186924 599768
rect 186780 584452 186832 584458
rect 186780 584394 186832 584400
rect 186792 526017 186820 584394
rect 186778 526008 186834 526017
rect 186778 525943 186834 525952
rect 186884 524385 186912 599762
rect 186976 599758 187004 608359
rect 186964 599752 187016 599758
rect 186964 599694 187016 599700
rect 186870 524376 186926 524385
rect 186870 524311 186926 524320
rect 186778 523288 186834 523297
rect 186778 523223 186834 523232
rect 186686 498264 186742 498273
rect 186686 498199 186742 498208
rect 186700 493270 186728 498199
rect 186688 493264 186740 493270
rect 186688 493206 186740 493212
rect 186792 489530 186820 523223
rect 186870 521520 186926 521529
rect 186870 521455 186926 521464
rect 186884 520305 186912 521455
rect 186870 520296 186926 520305
rect 186870 520231 186926 520240
rect 186884 494714 186912 520231
rect 186976 498273 187004 599694
rect 187068 599690 187096 610263
rect 187160 599962 187188 628623
rect 187252 600030 187280 631615
rect 187240 600024 187292 600030
rect 187240 599966 187292 599972
rect 187148 599956 187200 599962
rect 187148 599898 187200 599904
rect 187056 599684 187108 599690
rect 187056 599626 187108 599632
rect 187068 500313 187096 599626
rect 187160 518673 187188 599898
rect 187252 521665 187280 599966
rect 187344 599894 187372 637055
rect 187422 633312 187478 633321
rect 187422 633247 187478 633256
rect 187332 599888 187384 599894
rect 187332 599830 187384 599836
rect 187344 527105 187372 599830
rect 187330 527096 187386 527105
rect 187330 527031 187386 527040
rect 187344 525842 187372 527031
rect 187332 525836 187384 525842
rect 187332 525778 187384 525784
rect 187330 524376 187386 524385
rect 187330 524311 187386 524320
rect 187238 521656 187294 521665
rect 187238 521591 187294 521600
rect 187146 518664 187202 518673
rect 187146 518599 187202 518608
rect 187054 500304 187110 500313
rect 187054 500239 187110 500248
rect 186962 498264 187018 498273
rect 186962 498199 187018 498208
rect 186884 494686 187004 494714
rect 186872 493128 186924 493134
rect 186872 493070 186924 493076
rect 186780 489524 186832 489530
rect 186780 489466 186832 489472
rect 186792 488578 186820 489466
rect 186884 489462 186912 493070
rect 186976 489598 187004 494686
rect 187068 493406 187096 500239
rect 187056 493400 187108 493406
rect 187056 493342 187108 493348
rect 187056 493264 187108 493270
rect 187056 493206 187108 493212
rect 187068 489734 187096 493206
rect 187056 489728 187108 489734
rect 187056 489670 187108 489676
rect 186964 489592 187016 489598
rect 186964 489534 187016 489540
rect 186872 489456 186924 489462
rect 186872 489398 186924 489404
rect 186884 488782 186912 489398
rect 186872 488776 186924 488782
rect 186872 488718 186924 488724
rect 186780 488572 186832 488578
rect 186780 488514 186832 488520
rect 186976 449070 187004 489534
rect 187068 488646 187096 489670
rect 187160 489394 187188 518599
rect 187252 489802 187280 521591
rect 187240 489796 187292 489802
rect 187240 489738 187292 489744
rect 187148 489388 187200 489394
rect 187148 489330 187200 489336
rect 187056 488640 187108 488646
rect 187056 488582 187108 488588
rect 187160 449750 187188 489330
rect 187252 488714 187280 489738
rect 187344 489666 187372 524311
rect 187436 523297 187464 633247
rect 187514 630320 187570 630329
rect 187514 630255 187570 630264
rect 187422 523288 187478 523297
rect 187422 523223 187478 523232
rect 187528 521529 187556 630255
rect 187606 608696 187662 608705
rect 187606 608631 187662 608640
rect 187514 521520 187570 521529
rect 187514 521455 187570 521464
rect 187620 498681 187648 608631
rect 188620 596352 188672 596358
rect 188620 596294 188672 596300
rect 188528 596216 188580 596222
rect 188528 596158 188580 596164
rect 188344 581664 188396 581670
rect 188344 581606 188396 581612
rect 187700 525836 187752 525842
rect 187700 525778 187752 525784
rect 187606 498672 187662 498681
rect 187606 498607 187662 498616
rect 187712 489870 187740 525778
rect 187700 489864 187752 489870
rect 187700 489806 187752 489812
rect 187332 489660 187384 489666
rect 187332 489602 187384 489608
rect 187240 488708 187292 488714
rect 187240 488650 187292 488656
rect 187240 488572 187292 488578
rect 187240 488514 187292 488520
rect 187252 450770 187280 488514
rect 187240 450764 187292 450770
rect 187240 450706 187292 450712
rect 187344 450702 187372 489602
rect 187608 488776 187660 488782
rect 187608 488718 187660 488724
rect 187516 488708 187568 488714
rect 187516 488650 187568 488656
rect 187424 488640 187476 488646
rect 187424 488582 187476 488588
rect 187332 450696 187384 450702
rect 187332 450638 187384 450644
rect 187436 450634 187464 488582
rect 187528 450838 187556 488650
rect 187516 450832 187568 450838
rect 187516 450774 187568 450780
rect 187424 450628 187476 450634
rect 187424 450570 187476 450576
rect 187620 450566 187648 488718
rect 187712 486538 187740 489806
rect 187700 486532 187752 486538
rect 187700 486474 187752 486480
rect 187608 450560 187660 450566
rect 187608 450502 187660 450508
rect 187148 449744 187200 449750
rect 187148 449686 187200 449692
rect 188356 449546 188384 581606
rect 188434 526008 188490 526017
rect 188434 525943 188490 525952
rect 188448 450906 188476 525943
rect 188540 488442 188568 596158
rect 188632 488510 188660 596294
rect 188712 596284 188764 596290
rect 188712 596226 188764 596232
rect 188620 488504 188672 488510
rect 188620 488446 188672 488452
rect 188528 488436 188580 488442
rect 188528 488378 188580 488384
rect 188632 488238 188660 488446
rect 188620 488232 188672 488238
rect 188620 488174 188672 488180
rect 188724 488170 188752 596226
rect 188712 488164 188764 488170
rect 188712 488106 188764 488112
rect 188816 488102 188844 700266
rect 188804 488096 188856 488102
rect 188804 488038 188856 488044
rect 188436 450900 188488 450906
rect 188436 450842 188488 450848
rect 188344 449540 188396 449546
rect 188344 449482 188396 449488
rect 186964 449064 187016 449070
rect 186964 449006 187016 449012
rect 184204 448248 184256 448254
rect 184204 448190 184256 448196
rect 3976 448112 4028 448118
rect 3976 448054 4028 448060
rect 3792 447908 3844 447914
rect 3792 447850 3844 447856
rect 3240 447840 3292 447846
rect 3240 447782 3292 447788
rect 3700 446820 3752 446826
rect 3700 446762 3752 446768
rect 3424 446684 3476 446690
rect 3424 446626 3476 446632
rect 3240 445052 3292 445058
rect 3240 444994 3292 445000
rect 3252 423609 3280 444994
rect 3332 443080 3384 443086
rect 3332 443022 3384 443028
rect 3238 423600 3294 423609
rect 3238 423535 3294 423544
rect 2780 410984 2832 410990
rect 2780 410926 2832 410932
rect 2792 410553 2820 410926
rect 2778 410544 2834 410553
rect 2778 410479 2834 410488
rect 3344 397497 3372 443022
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3148 267708 3200 267714
rect 3148 267650 3200 267656
rect 3160 267209 3188 267650
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3056 215280 3108 215286
rect 3056 215222 3108 215228
rect 3068 214985 3096 215222
rect 3054 214976 3110 214985
rect 3054 214911 3110 214920
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3436 84697 3464 446626
rect 3514 446448 3570 446457
rect 3514 446383 3570 446392
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3528 45529 3556 446383
rect 3608 443012 3660 443018
rect 3608 442954 3660 442960
rect 3620 136785 3648 442954
rect 3712 188873 3740 446762
rect 4988 446616 5040 446622
rect 4988 446558 5040 446564
rect 4896 446140 4948 446146
rect 4896 446082 4948 446088
rect 3884 446072 3936 446078
rect 3884 446014 3936 446020
rect 3792 445868 3844 445874
rect 3792 445810 3844 445816
rect 3804 201929 3832 445810
rect 3896 241097 3924 446014
rect 4804 445936 4856 445942
rect 4804 445878 4856 445884
rect 3976 445120 4028 445126
rect 3976 445062 4028 445068
rect 3988 254153 4016 445062
rect 4068 443148 4120 443154
rect 4068 443090 4120 443096
rect 4080 345409 4108 443090
rect 4160 393984 4212 393990
rect 4160 393926 4212 393932
rect 4066 345400 4122 345409
rect 4066 345335 4122 345344
rect 3974 254144 4030 254153
rect 3974 254079 4030 254088
rect 3882 241088 3938 241097
rect 3882 241023 3938 241032
rect 3790 201920 3846 201929
rect 3790 201855 3846 201864
rect 3698 188864 3754 188873
rect 3698 188799 3754 188808
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 393926
rect 4816 97782 4844 445878
rect 4908 358494 4936 446082
rect 5000 410990 5028 446558
rect 188908 446486 188936 700402
rect 218992 700398 219020 703520
rect 188988 700392 189040 700398
rect 188988 700334 189040 700340
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 188896 446480 188948 446486
rect 188896 446422 188948 446428
rect 189000 446418 189028 700334
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 207846 597544 207902 597553
rect 207846 597479 207902 597488
rect 208950 597544 209006 597553
rect 208950 597479 209006 597488
rect 209962 597544 210018 597553
rect 209962 597479 210018 597488
rect 211158 597544 211214 597553
rect 211158 597479 211214 597488
rect 212354 597544 212410 597553
rect 212354 597479 212410 597488
rect 213826 597544 213882 597553
rect 213826 597479 213882 597488
rect 214838 597544 214894 597553
rect 214838 597479 214894 597488
rect 215298 597544 215354 597553
rect 215298 597479 215354 597488
rect 215758 597544 215814 597553
rect 215758 597479 215814 597488
rect 226246 597544 226302 597553
rect 226246 597479 226302 597488
rect 235906 597544 235962 597553
rect 235906 597479 235962 597488
rect 245566 597544 245622 597553
rect 245566 597479 245622 597488
rect 251086 597544 251142 597553
rect 251086 597479 251142 597488
rect 204350 597136 204406 597145
rect 204350 597071 204406 597080
rect 202878 596456 202934 596465
rect 202878 596391 202934 596400
rect 202892 596358 202920 596391
rect 202880 596352 202932 596358
rect 202880 596294 202932 596300
rect 204258 596320 204314 596329
rect 204364 596290 204392 597071
rect 207860 596834 207888 597479
rect 208964 597106 208992 597479
rect 209976 597174 210004 597479
rect 209964 597168 210016 597174
rect 209964 597110 210016 597116
rect 211068 597168 211120 597174
rect 211068 597110 211120 597116
rect 208952 597100 209004 597106
rect 208952 597042 209004 597048
rect 207848 596828 207900 596834
rect 207848 596770 207900 596776
rect 204258 596255 204314 596264
rect 204352 596284 204404 596290
rect 204272 596222 204300 596255
rect 204352 596226 204404 596232
rect 207860 596222 207888 596770
rect 208964 596358 208992 597042
rect 208952 596352 209004 596358
rect 208952 596294 209004 596300
rect 211080 596290 211108 597110
rect 211172 597038 211200 597479
rect 212368 597310 212396 597479
rect 212356 597304 212408 597310
rect 212356 597246 212408 597252
rect 211160 597032 211212 597038
rect 211160 596974 211212 596980
rect 212368 596426 212396 597246
rect 213840 597038 213868 597479
rect 214852 597242 214880 597479
rect 214840 597236 214892 597242
rect 214840 597178 214892 597184
rect 212448 597032 212500 597038
rect 212448 596974 212500 596980
rect 213828 597032 213880 597038
rect 213828 596974 213880 596980
rect 212460 596834 212488 596974
rect 213840 596902 213868 596974
rect 214852 596902 214880 597178
rect 213828 596896 213880 596902
rect 213828 596838 213880 596844
rect 214840 596896 214892 596902
rect 214840 596838 214892 596844
rect 212448 596828 212500 596834
rect 212448 596770 212500 596776
rect 212356 596420 212408 596426
rect 212356 596362 212408 596368
rect 211068 596284 211120 596290
rect 211068 596226 211120 596232
rect 204260 596216 204312 596222
rect 204260 596158 204312 596164
rect 207848 596216 207900 596222
rect 207848 596158 207900 596164
rect 215312 580378 215340 597479
rect 215772 596970 215800 597479
rect 215760 596964 215812 596970
rect 215760 596906 215812 596912
rect 219438 596320 219494 596329
rect 219438 596255 219494 596264
rect 190000 580372 190052 580378
rect 190000 580314 190052 580320
rect 215300 580372 215352 580378
rect 215300 580314 215352 580320
rect 189908 580304 189960 580310
rect 189908 580246 189960 580252
rect 189078 498672 189134 498681
rect 189078 498607 189134 498616
rect 189092 450974 189120 498607
rect 189080 450968 189132 450974
rect 189080 450910 189132 450916
rect 189920 449682 189948 580246
rect 189908 449676 189960 449682
rect 189908 449618 189960 449624
rect 190012 449614 190040 580314
rect 219452 580310 219480 596255
rect 226260 581670 226288 597479
rect 231766 597272 231822 597281
rect 231766 597207 231822 597216
rect 226248 581664 226300 581670
rect 226248 581606 226300 581612
rect 231780 580310 231808 597207
rect 235920 580378 235948 597479
rect 241426 596864 241482 596873
rect 241426 596799 241482 596808
rect 241440 580446 241468 596799
rect 245580 580514 245608 597479
rect 251100 580582 251128 597479
rect 280988 597372 281040 597378
rect 280988 597314 281040 597320
rect 251088 580576 251140 580582
rect 251088 580518 251140 580524
rect 245568 580508 245620 580514
rect 245568 580450 245620 580456
rect 241428 580440 241480 580446
rect 241428 580382 241480 580388
rect 235908 580372 235960 580378
rect 235908 580314 235960 580320
rect 219440 580304 219492 580310
rect 219440 580246 219492 580252
rect 231768 580304 231820 580310
rect 231768 580246 231820 580252
rect 253664 489252 253716 489258
rect 253664 489194 253716 489200
rect 218060 489184 218112 489190
rect 218060 489126 218112 489132
rect 204718 488472 204774 488481
rect 204718 488407 204720 488416
rect 204772 488407 204774 488416
rect 214838 488472 214894 488481
rect 214838 488407 214894 488416
rect 204720 488378 204772 488384
rect 202880 488232 202932 488238
rect 202878 488200 202880 488209
rect 202932 488200 202934 488209
rect 202878 488135 202934 488144
rect 204732 487286 204760 488378
rect 211158 488336 211214 488345
rect 211158 488271 211214 488280
rect 213734 488336 213790 488345
rect 213734 488271 213790 488280
rect 204904 488164 204956 488170
rect 204904 488106 204956 488112
rect 204720 487280 204772 487286
rect 203522 487248 203578 487257
rect 204916 487257 204944 488106
rect 208858 487928 208914 487937
rect 208858 487863 208914 487872
rect 207664 487484 207716 487490
rect 207664 487426 207716 487432
rect 207676 487257 207704 487426
rect 208872 487354 208900 487863
rect 211172 487830 211200 488271
rect 213748 487898 213776 488271
rect 214852 487966 214880 488407
rect 215758 488336 215814 488345
rect 215758 488271 215814 488280
rect 215772 488034 215800 488271
rect 215760 488028 215812 488034
rect 215760 487970 215812 487976
rect 214840 487960 214892 487966
rect 214840 487902 214892 487908
rect 213736 487892 213788 487898
rect 213736 487834 213788 487840
rect 211160 487824 211212 487830
rect 211160 487766 211212 487772
rect 212448 487824 212500 487830
rect 212448 487766 212500 487772
rect 212354 487520 212410 487529
rect 212354 487455 212410 487464
rect 212368 487422 212396 487455
rect 212460 487422 212488 487766
rect 212356 487416 212408 487422
rect 212356 487358 212408 487364
rect 212448 487416 212500 487422
rect 212448 487358 212500 487364
rect 208860 487348 208912 487354
rect 208860 487290 208912 487296
rect 204720 487222 204772 487228
rect 204902 487248 204958 487257
rect 203522 487183 203578 487192
rect 204902 487183 204958 487192
rect 207662 487248 207718 487257
rect 207662 487183 207718 487192
rect 203536 459474 203564 487183
rect 203524 459468 203576 459474
rect 203524 459410 203576 459416
rect 190000 449608 190052 449614
rect 190000 449550 190052 449556
rect 204916 449138 204944 487183
rect 207676 460902 207704 487183
rect 208872 486606 208900 487290
rect 210422 487248 210478 487257
rect 210422 487183 210424 487192
rect 210476 487183 210478 487192
rect 210424 487154 210476 487160
rect 208860 486600 208912 486606
rect 208860 486542 208912 486548
rect 207664 460896 207716 460902
rect 207664 460838 207716 460844
rect 210436 459542 210464 487154
rect 212368 483750 212396 487358
rect 213748 487354 213776 487834
rect 214852 487490 214880 487902
rect 214840 487484 214892 487490
rect 214840 487426 214892 487432
rect 213736 487348 213788 487354
rect 213736 487290 213788 487296
rect 215772 487218 215800 487970
rect 216586 487248 216642 487257
rect 215760 487212 215812 487218
rect 216586 487183 216642 487192
rect 215760 487154 215812 487160
rect 212356 483744 212408 483750
rect 212356 483686 212408 483692
rect 215300 480956 215352 480962
rect 215300 480898 215352 480904
rect 214012 470620 214064 470626
rect 214012 470562 214064 470568
rect 210424 459536 210476 459542
rect 210424 459478 210476 459484
rect 204904 449132 204956 449138
rect 204904 449074 204956 449080
rect 213184 447772 213236 447778
rect 213184 447714 213236 447720
rect 211712 447704 211764 447710
rect 211712 447646 211764 447652
rect 211158 447264 211214 447273
rect 211158 447199 211214 447208
rect 188988 446412 189040 446418
rect 188988 446354 189040 446360
rect 210422 446312 210478 446321
rect 210422 446247 210478 446256
rect 209134 446176 209190 446185
rect 209134 446111 209190 446120
rect 79322 446040 79378 446049
rect 79322 445975 79378 445984
rect 4988 410984 5040 410990
rect 4988 410926 5040 410932
rect 25502 397488 25558 397497
rect 25502 397423 25558 397432
rect 13818 392592 13874 392601
rect 13818 392527 13874 392536
rect 4896 358488 4948 358494
rect 4896 358430 4948 358436
rect 5540 352572 5592 352578
rect 5540 352514 5592 352520
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 5552 16574 5580 352514
rect 9680 177336 9732 177342
rect 9680 177278 9732 177284
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 3608 13116 3660 13122
rect 3608 13058 3660 13064
rect 1674 9072 1730 9081
rect 1674 9007 1730 9016
rect 570 8936 626 8945
rect 570 8871 626 8880
rect 584 480 612 8871
rect 1688 480 1716 9007
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 480 2912 8910
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 13058
rect 5276 480 5304 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 480 7696 8978
rect 8772 480 8800 13126
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 177278
rect 13832 16574 13860 392527
rect 23480 338768 23532 338774
rect 23480 338710 23532 338716
rect 23492 16574 23520 338710
rect 24860 333260 24912 333266
rect 24860 333202 24912 333208
rect 24872 16574 24900 333202
rect 13832 16546 14320 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 11152 10328 11204 10334
rect 11152 10270 11204 10276
rect 11164 480 11192 10270
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 480 13584 3470
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 480 15976 12038
rect 17038 11656 17094 11665
rect 17038 11591 17094 11600
rect 17052 480 17080 11591
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 14418
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19444 480 19472 4762
rect 20628 3256 20680 3262
rect 20628 3198 20680 3204
rect 20640 480 20668 3198
rect 21836 480 21864 11698
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 14486
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3262 25544 397423
rect 77300 396908 77352 396914
rect 77300 396850 77352 396856
rect 46940 396840 46992 396846
rect 46940 396782 46992 396788
rect 40040 396772 40092 396778
rect 40040 396714 40092 396720
rect 30380 395412 30432 395418
rect 30380 395354 30432 395360
rect 27620 395344 27672 395350
rect 27620 395286 27672 395292
rect 27710 395312 27766 395321
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 25504 3256 25556 3262
rect 25504 3198 25556 3204
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 11766
rect 27632 6914 27660 395286
rect 27710 395247 27766 395256
rect 27724 16574 27752 395247
rect 30392 16574 30420 395354
rect 37280 355360 37332 355366
rect 37280 355302 37332 355308
rect 31760 169040 31812 169046
rect 31760 168982 31812 168988
rect 31772 16574 31800 168982
rect 37292 16574 37320 355302
rect 38660 181484 38712 181490
rect 38660 181426 38712 181432
rect 38672 16574 38700 181426
rect 40052 16574 40080 396714
rect 45558 395448 45614 395457
rect 45558 395383 45614 395392
rect 42800 355428 42852 355434
rect 42800 355370 42852 355376
rect 41420 178696 41472 178702
rect 41420 178638 41472 178644
rect 41432 16574 41460 178638
rect 27724 16546 28488 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30102 11792 30158 11801
rect 30102 11727 30158 11736
rect 30116 480 30144 11727
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 34520 14612 34572 14618
rect 34520 14554 34572 14560
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 33612 480 33640 11834
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 14554
rect 36004 480 36032 15846
rect 36728 11960 36780 11966
rect 36728 11902 36780 11908
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 11902
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 355370
rect 45572 16574 45600 395383
rect 46952 16574 46980 396782
rect 64878 396672 64934 396681
rect 64878 396607 64934 396616
rect 52460 395480 52512 395486
rect 52460 395422 52512 395428
rect 52472 16574 52500 395422
rect 60740 354136 60792 354142
rect 60740 354078 60792 354084
rect 56600 354000 56652 354006
rect 56600 353942 56652 353948
rect 56612 16574 56640 353942
rect 60752 16574 60780 354078
rect 62120 354068 62172 354074
rect 62120 354010 62172 354016
rect 62132 16574 62160 354010
rect 63498 177304 63554 177313
rect 63498 177239 63554 177248
rect 63512 16574 63540 177239
rect 64892 16574 64920 396607
rect 67638 395584 67694 395593
rect 67638 395519 67694 395528
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 52472 16546 53328 16574
rect 56612 16546 56824 16574
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 44180 14680 44232 14686
rect 44180 14622 44232 14628
rect 44192 3466 44220 14622
rect 44272 12028 44324 12034
rect 44272 11970 44324 11976
rect 44180 3460 44232 3466
rect 44180 3402 44232 3408
rect 44284 480 44312 11970
rect 45100 3460 45152 3466
rect 45100 3402 45152 3408
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3402
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 50158 14512 50214 14521
rect 50158 14447 50214 14456
rect 48502 11928 48558 11937
rect 48502 11863 48558 11872
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 11863
rect 50172 480 50200 14447
rect 51354 7576 51410 7585
rect 51354 7511 51410 7520
rect 51368 480 51396 7511
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 52564 480 52592 3402
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 56048 13252 56100 13258
rect 56048 13194 56100 13200
rect 54944 7608 54996 7614
rect 54944 7550 54996 7556
rect 54956 480 54984 7550
rect 56060 480 56088 13194
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 59360 13320 59412 13326
rect 59360 13262 59412 13268
rect 58440 9104 58492 9110
rect 58440 9046 58492 9052
rect 58452 480 58480 9046
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13262
rect 60844 480 60872 16546
rect 62028 9172 62080 9178
rect 62028 9114 62080 9120
rect 62040 480 62068 9114
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66718 13016 66774 13025
rect 66718 12951 66774 12960
rect 66732 480 66760 12951
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 395519
rect 69020 394052 69072 394058
rect 69020 393994 69072 394000
rect 69032 16574 69060 393994
rect 70400 354204 70452 354210
rect 70400 354146 70452 354152
rect 70412 16574 70440 354146
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 69124 480 69152 16546
rect 69848 13388 69900 13394
rect 69848 13330 69900 13336
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 13330
rect 71516 480 71544 16546
rect 75000 14748 75052 14754
rect 75000 14690 75052 14696
rect 73344 13456 73396 13462
rect 73344 13398 73396 13404
rect 72608 9240 72660 9246
rect 72608 9182 72660 9188
rect 72620 480 72648 9182
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 13398
rect 75012 480 75040 14690
rect 76196 9308 76248 9314
rect 76196 9250 76248 9256
rect 76208 480 76236 9250
rect 77312 3398 77340 396850
rect 79336 59362 79364 445975
rect 196716 445324 196768 445330
rect 196716 445266 196768 445272
rect 98644 445256 98696 445262
rect 98644 445198 98696 445204
rect 98656 372570 98684 445198
rect 196624 444576 196676 444582
rect 196624 444518 196676 444524
rect 192484 443216 192536 443222
rect 192484 443158 192536 443164
rect 189080 398336 189132 398342
rect 188342 398304 188398 398313
rect 171140 398268 171192 398274
rect 189080 398278 189132 398284
rect 188342 398239 188398 398248
rect 171140 398210 171192 398216
rect 164240 398200 164292 398206
rect 164240 398142 164292 398148
rect 125600 398132 125652 398138
rect 125600 398074 125652 398080
rect 100758 396808 100814 396817
rect 100758 396743 100814 396752
rect 98644 372564 98696 372570
rect 98644 372506 98696 372512
rect 92480 355496 92532 355502
rect 92480 355438 92532 355444
rect 88340 354408 88392 354414
rect 88340 354350 88392 354356
rect 86960 354272 87012 354278
rect 86960 354214 87012 354220
rect 84198 353968 84254 353977
rect 84198 353903 84254 353912
rect 79324 59356 79376 59362
rect 79324 59298 79376 59304
rect 80888 13592 80940 13598
rect 80888 13534 80940 13540
rect 77392 13524 77444 13530
rect 77392 13466 77444 13472
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 13466
rect 79692 9376 79744 9382
rect 79692 9318 79744 9324
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 79704 480 79732 9318
rect 80900 480 80928 13534
rect 83278 10296 83334 10305
rect 83278 10231 83334 10240
rect 82084 3800 82136 3806
rect 82084 3742 82136 3748
rect 82096 480 82124 3742
rect 83292 480 83320 10231
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 353903
rect 85580 351212 85632 351218
rect 85580 351154 85632 351160
rect 85592 16574 85620 351154
rect 86972 16574 87000 354214
rect 88352 16574 88380 354350
rect 91100 354340 91152 354346
rect 91100 354282 91152 354288
rect 91112 16574 91140 354282
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 88932 16574
rect 91112 16546 91600 16574
rect 85684 480 85712 16546
rect 86406 10432 86462 10441
rect 86406 10367 86462 10376
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 10367
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 88246 9208 88302 9217
rect 88246 9143 88302 9152
rect 88260 3602 88288 9143
rect 88248 3596 88300 3602
rect 88248 3538 88300 3544
rect 88904 3482 88932 16546
rect 88982 13152 89038 13161
rect 88982 13087 89038 13096
rect 88996 3602 89024 13087
rect 89904 10396 89956 10402
rect 89904 10338 89956 10344
rect 88984 3596 89036 3602
rect 88984 3538 89036 3544
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 10338
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 355438
rect 95240 83496 95292 83502
rect 95240 83438 95292 83444
rect 95252 16574 95280 83438
rect 95252 16546 95832 16574
rect 93952 10464 94004 10470
rect 93952 10406 94004 10412
rect 93964 480 93992 10406
rect 95148 4004 95200 4010
rect 95148 3946 95200 3952
rect 95160 480 95188 3946
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 99838 15872 99894 15881
rect 99838 15807 99894 15816
rect 98184 14816 98236 14822
rect 98184 14758 98236 14764
rect 97448 10532 97500 10538
rect 97448 10474 97500 10480
rect 97460 480 97488 10474
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 14758
rect 99852 480 99880 15807
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 396743
rect 118698 395720 118754 395729
rect 118698 395655 118754 395664
rect 115940 395548 115992 395554
rect 115940 395490 115992 395496
rect 109040 392624 109092 392630
rect 109040 392566 109092 392572
rect 106280 363656 106332 363662
rect 106280 363598 106332 363604
rect 102138 354104 102194 354113
rect 102138 354039 102194 354048
rect 102152 6914 102180 354039
rect 102232 180124 102284 180130
rect 102232 180066 102284 180072
rect 102244 16574 102272 180066
rect 106292 16574 106320 363598
rect 102244 16546 103376 16574
rect 106292 16546 106504 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 105728 14884 105780 14890
rect 105728 14826 105780 14832
rect 104072 10600 104124 10606
rect 104072 10542 104124 10548
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 10542
rect 105740 480 105768 14826
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 10668 108172 10674
rect 108120 10610 108172 10616
rect 108132 480 108160 10610
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 392566
rect 110420 340196 110472 340202
rect 110420 340138 110472 340144
rect 110432 16574 110460 340138
rect 115952 16574 115980 395490
rect 117320 86284 117372 86290
rect 117320 86226 117372 86232
rect 110432 16546 110552 16574
rect 115952 16546 116440 16574
rect 110524 480 110552 16546
rect 114008 15972 114060 15978
rect 114008 15914 114060 15920
rect 111616 10736 111668 10742
rect 111616 10678 111668 10684
rect 111628 480 111656 10678
rect 112812 3868 112864 3874
rect 112812 3810 112864 3816
rect 112824 480 112852 3810
rect 114020 480 114048 15914
rect 115204 3936 115256 3942
rect 115204 3878 115256 3884
rect 115216 480 115244 3878
rect 116412 480 116440 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 86226
rect 118712 3534 118740 395655
rect 120078 177440 120134 177449
rect 120078 177375 120134 177384
rect 124220 177404 124272 177410
rect 120092 16574 120120 177375
rect 124220 177346 124272 177352
rect 124232 16574 124260 177346
rect 120092 16546 120672 16574
rect 124232 16546 124720 16574
rect 118792 3732 118844 3738
rect 118792 3674 118844 3680
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 118804 480 118832 3674
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 119908 480 119936 3470
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 123024 14952 123076 14958
rect 123024 14894 123076 14900
rect 122286 12064 122342 12073
rect 122286 11999 122342 12008
rect 122300 480 122328 11999
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 14894
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 398074
rect 155960 397112 156012 397118
rect 155960 397054 156012 397060
rect 144920 397044 144972 397050
rect 144920 396986 144972 396992
rect 131120 396976 131172 396982
rect 131120 396918 131172 396924
rect 129740 394120 129792 394126
rect 129740 394062 129792 394068
rect 129752 16574 129780 394062
rect 131132 16574 131160 396918
rect 139398 394088 139454 394097
rect 139398 394023 139454 394032
rect 135258 393952 135314 393961
rect 135258 393887 135314 393896
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 128176 6180 128228 6186
rect 128176 6122 128228 6128
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 6122
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 129384 480 129412 3538
rect 130580 480 130608 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 134156 6248 134208 6254
rect 134156 6190 134208 6196
rect 132960 4888 133012 4894
rect 132960 4830 133012 4836
rect 132972 480 133000 4830
rect 134168 480 134196 6190
rect 135272 3398 135300 393887
rect 139412 16574 139440 394023
rect 140780 177472 140832 177478
rect 140780 177414 140832 177420
rect 140792 16574 140820 177414
rect 144932 16574 144960 396986
rect 149704 395616 149756 395622
rect 149704 395558 149756 395564
rect 149060 46232 149112 46238
rect 149060 46174 149112 46180
rect 149072 16574 149100 46174
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 144932 16546 145512 16574
rect 149072 16546 149560 16574
rect 138662 14648 138718 14657
rect 138662 14583 138718 14592
rect 137650 7712 137706 7721
rect 137650 7647 137706 7656
rect 135352 3664 135404 3670
rect 135352 3606 135404 3612
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 135364 1714 135392 3606
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 135272 1686 135392 1714
rect 135272 480 135300 1686
rect 136468 480 136496 3334
rect 137664 480 137692 7647
rect 138676 3806 138704 14583
rect 138846 7848 138902 7857
rect 138846 7783 138902 7792
rect 138664 3800 138716 3806
rect 138664 3742 138716 3748
rect 138860 480 138888 7783
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 144736 7744 144788 7750
rect 144736 7686 144788 7692
rect 142436 7676 142488 7682
rect 142436 7618 142488 7624
rect 142448 480 142476 7618
rect 143540 4956 143592 4962
rect 143540 4898 143592 4904
rect 143552 480 143580 4898
rect 144748 480 144776 7686
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 148324 7812 148376 7818
rect 148324 7754 148376 7760
rect 147128 5160 147180 5166
rect 147128 5102 147180 5108
rect 147140 480 147168 5102
rect 148336 480 148364 7754
rect 149532 480 149560 16546
rect 149716 4010 149744 395558
rect 153198 394224 153254 394233
rect 153198 394159 153254 394168
rect 151818 392728 151874 392737
rect 151818 392663 151874 392672
rect 150624 5228 150676 5234
rect 150624 5170 150676 5176
rect 149704 4004 149756 4010
rect 149704 3946 149756 3952
rect 150636 480 150664 5170
rect 151832 3806 151860 392663
rect 153212 16574 153240 394159
rect 154580 177540 154632 177546
rect 154580 177482 154632 177488
rect 154592 16574 154620 177482
rect 155972 16574 156000 397054
rect 160100 392692 160152 392698
rect 160100 392634 160152 392640
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 151912 7880 151964 7886
rect 151912 7822 151964 7828
rect 151820 3800 151872 3806
rect 151820 3742 151872 3748
rect 151924 3482 151952 7822
rect 153016 3800 153068 3806
rect 153016 3742 153068 3748
rect 151832 3454 151952 3482
rect 151832 480 151860 3454
rect 153028 480 153056 3742
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 160112 11694 160140 392634
rect 160192 352640 160244 352646
rect 160192 352582 160244 352588
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 158904 7948 158956 7954
rect 158904 7890 158956 7896
rect 157800 5160 157852 5166
rect 157800 5102 157852 5108
rect 157812 480 157840 5102
rect 158916 480 158944 7890
rect 160204 6914 160232 352582
rect 162860 46300 162912 46306
rect 162860 46242 162912 46248
rect 162872 16574 162900 46242
rect 164252 16574 164280 398142
rect 169024 354476 169076 354482
rect 169024 354418 169076 354424
rect 167000 177608 167052 177614
rect 167000 177550 167052 177556
rect 167012 16574 167040 177550
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 167012 16546 167224 16574
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11630
rect 162492 5228 162544 5234
rect 162492 5170 162544 5176
rect 162504 480 162532 5170
rect 163700 480 163728 16546
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166080 5296 166132 5302
rect 166080 5238 166132 5244
rect 166092 480 166120 5238
rect 167196 480 167224 16546
rect 169036 3874 169064 354418
rect 171152 16574 171180 398210
rect 178682 398168 178738 398177
rect 178682 398103 178738 398112
rect 178040 394188 178092 394194
rect 178040 394130 178092 394136
rect 176660 178764 176712 178770
rect 176660 178706 176712 178712
rect 173898 177576 173954 177585
rect 173898 177511 173954 177520
rect 171152 16546 171732 16574
rect 170310 16008 170366 16017
rect 170310 15943 170366 15952
rect 169576 6316 169628 6322
rect 169576 6258 169628 6264
rect 169024 3868 169076 3874
rect 169024 3810 169076 3816
rect 168380 3800 168432 3806
rect 168380 3742 168432 3748
rect 168392 480 168420 3742
rect 169588 480 169616 6258
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 15943
rect 171704 3482 171732 16546
rect 171784 10804 171836 10810
rect 171784 10746 171836 10752
rect 171796 3942 171824 10746
rect 173162 6216 173218 6225
rect 173162 6151 173218 6160
rect 171784 3936 171836 3942
rect 171784 3878 171836 3884
rect 171704 3454 172008 3482
rect 171980 480 172008 3454
rect 173176 480 173204 6151
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 177511
rect 176672 3466 176700 178706
rect 178052 16574 178080 394130
rect 178052 16546 178632 16574
rect 176752 6384 176804 6390
rect 176752 6326 176804 6332
rect 176660 3460 176712 3466
rect 176660 3402 176712 3408
rect 175462 3360 175518 3369
rect 175462 3295 175518 3304
rect 175476 480 175504 3295
rect 176764 3210 176792 6326
rect 177856 3460 177908 3466
rect 177856 3402 177908 3408
rect 176672 3182 176792 3210
rect 176672 480 176700 3182
rect 177868 480 177896 3402
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 12102 178724 398103
rect 180800 352708 180852 352714
rect 180800 352650 180852 352656
rect 180812 16574 180840 352650
rect 187698 178664 187754 178673
rect 187698 178599 187754 178608
rect 180812 16546 181024 16574
rect 178684 12096 178736 12102
rect 178684 12038 178736 12044
rect 178776 12096 178828 12102
rect 178776 12038 178828 12044
rect 178788 3398 178816 12038
rect 180248 6452 180300 6458
rect 180248 6394 180300 6400
rect 178776 3392 178828 3398
rect 178776 3334 178828 3340
rect 180260 480 180288 6394
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 185582 10568 185638 10577
rect 185582 10503 185638 10512
rect 183744 6520 183796 6526
rect 183744 6462 183796 6468
rect 182548 3460 182600 3466
rect 182548 3402 182600 3408
rect 182560 480 182588 3402
rect 183756 480 183784 6462
rect 184940 3868 184992 3874
rect 184940 3810 184992 3816
rect 184952 480 184980 3810
rect 185596 3738 185624 10503
rect 187712 6914 187740 178599
rect 188356 10334 188384 398239
rect 189092 16574 189120 398278
rect 191838 352608 191894 352617
rect 191838 352543 191894 352552
rect 190458 46200 190514 46209
rect 190458 46135 190514 46144
rect 189092 16546 189304 16574
rect 188344 10328 188396 10334
rect 188344 10270 188396 10276
rect 187712 6886 188568 6914
rect 187332 6588 187384 6594
rect 187332 6530 187384 6536
rect 186136 3936 186188 3942
rect 186136 3878 186188 3884
rect 185584 3732 185636 3738
rect 185584 3674 185636 3680
rect 186148 480 186176 3878
rect 187344 480 187372 6530
rect 188540 480 188568 6886
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 46135
rect 191852 16574 191880 352543
rect 192496 150414 192524 443158
rect 194600 397180 194652 397186
rect 194600 397122 194652 397128
rect 193220 394256 193272 394262
rect 193220 394198 193272 394204
rect 192484 150408 192536 150414
rect 192484 150350 192536 150356
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 394198
rect 194612 16574 194640 397122
rect 196636 164218 196664 444518
rect 196728 267714 196756 445266
rect 199568 445188 199620 445194
rect 199568 445130 199620 445136
rect 199476 444916 199528 444922
rect 199476 444858 199528 444864
rect 199384 444848 199436 444854
rect 199384 444790 199436 444796
rect 198004 443284 198056 443290
rect 198004 443226 198056 443232
rect 196716 267708 196768 267714
rect 196716 267650 196768 267656
rect 196624 164212 196676 164218
rect 196624 164154 196676 164160
rect 198016 33114 198044 443226
rect 198740 352776 198792 352782
rect 198740 352718 198792 352724
rect 198004 33108 198056 33114
rect 198004 33050 198056 33056
rect 194612 16546 195192 16574
rect 194414 6352 194470 6361
rect 194414 6287 194470 6296
rect 194428 480 194456 6287
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 197912 8016 197964 8022
rect 197912 7958 197964 7964
rect 196808 5364 196860 5370
rect 196808 5306 196860 5312
rect 196820 480 196848 5306
rect 197924 480 197952 7958
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 352718
rect 199396 111790 199424 444790
rect 199488 215286 199516 444858
rect 199580 320142 199608 445130
rect 200856 444440 200908 444446
rect 200856 444382 200908 444388
rect 200764 443352 200816 443358
rect 200764 443294 200816 443300
rect 199568 320136 199620 320142
rect 199568 320078 199620 320084
rect 199476 215280 199528 215286
rect 199476 215222 199528 215228
rect 199384 111784 199436 111790
rect 199384 111726 199436 111732
rect 200776 20670 200804 443294
rect 200868 71738 200896 444382
rect 209148 443972 209176 446111
rect 210054 444952 210110 444961
rect 210054 444887 210110 444896
rect 209686 444816 209742 444825
rect 209686 444751 209742 444760
rect 209502 444136 209558 444145
rect 209332 444060 209452 444088
rect 209502 444071 209558 444080
rect 209332 443972 209360 444060
rect 209424 443873 209452 444060
rect 209516 443972 209544 444071
rect 209700 443972 209728 444751
rect 209884 444060 210004 444088
rect 209884 443972 209912 444060
rect 209410 443864 209466 443873
rect 209410 443799 209466 443808
rect 209976 443601 210004 444060
rect 210068 443972 210096 444887
rect 210238 444680 210294 444689
rect 210238 444615 210294 444624
rect 210252 443972 210280 444615
rect 210436 443972 210464 446247
rect 210790 444544 210846 444553
rect 210790 444479 210846 444488
rect 210606 444136 210662 444145
rect 210606 444071 210662 444080
rect 210620 443972 210648 444071
rect 210804 443972 210832 444479
rect 210988 444060 211108 444088
rect 210988 443972 211016 444060
rect 209962 443592 210018 443601
rect 209962 443527 210018 443536
rect 211080 443465 211108 444060
rect 211172 443972 211200 447199
rect 211528 445392 211580 445398
rect 211528 445334 211580 445340
rect 211344 444712 211396 444718
rect 211344 444654 211396 444660
rect 211356 443972 211384 444654
rect 211540 443972 211568 445334
rect 211724 443972 211752 447646
rect 212816 447636 212868 447642
rect 212816 447578 212868 447584
rect 212632 447568 212684 447574
rect 212632 447510 212684 447516
rect 212264 447500 212316 447506
rect 212264 447442 212316 447448
rect 212080 446344 212132 446350
rect 212080 446286 212132 446292
rect 211896 444780 211948 444786
rect 211896 444722 211948 444728
rect 211908 443972 211936 444722
rect 212092 443972 212120 446286
rect 212276 443972 212304 447442
rect 212368 444060 212488 444088
rect 212368 443465 212396 444060
rect 212460 443972 212488 444060
rect 212644 443972 212672 447510
rect 212828 443972 212856 447578
rect 213000 444984 213052 444990
rect 213000 444926 213052 444932
rect 213012 443972 213040 444926
rect 213196 443972 213224 447714
rect 214024 447370 214052 470562
rect 214196 460216 214248 460222
rect 214196 460158 214248 460164
rect 214012 447364 214064 447370
rect 214012 447306 214064 447312
rect 214208 447302 214236 460158
rect 214288 455524 214340 455530
rect 214288 455466 214340 455472
rect 214196 447296 214248 447302
rect 214196 447238 214248 447244
rect 213736 447160 213788 447166
rect 213736 447102 213788 447108
rect 213368 446276 213420 446282
rect 213368 446218 213420 446224
rect 213380 443972 213408 446218
rect 213564 444060 213684 444088
rect 213564 443972 213592 444060
rect 213656 443465 213684 444060
rect 213748 443972 213776 447102
rect 214104 446208 214156 446214
rect 214104 446150 214156 446156
rect 213920 444508 213972 444514
rect 213920 444450 213972 444456
rect 213932 443972 213960 444450
rect 214116 443972 214144 446150
rect 214300 443972 214328 455466
rect 214472 455456 214524 455462
rect 214472 455398 214524 455404
rect 214484 443972 214512 455398
rect 214656 453348 214708 453354
rect 214656 453290 214708 453296
rect 214668 443972 214696 453290
rect 214840 451308 214892 451314
rect 214840 451250 214892 451256
rect 214852 443972 214880 451250
rect 215024 447364 215076 447370
rect 215024 447306 215076 447312
rect 215036 443972 215064 447306
rect 215208 447296 215260 447302
rect 215208 447238 215260 447244
rect 215220 443972 215248 447238
rect 215312 447234 215340 480898
rect 215484 479528 215536 479534
rect 215484 479470 215536 479476
rect 215392 472660 215444 472666
rect 215392 472602 215444 472608
rect 215300 447228 215352 447234
rect 215300 447170 215352 447176
rect 215404 443972 215432 472602
rect 215496 460934 215524 479470
rect 215668 474020 215720 474026
rect 215668 473962 215720 473968
rect 215496 460906 215616 460934
rect 215588 443972 215616 460906
rect 215680 447370 215708 473962
rect 216600 472802 216628 487183
rect 216772 486464 216824 486470
rect 216772 486406 216824 486412
rect 216680 482316 216732 482322
rect 216680 482258 216732 482264
rect 216588 472796 216640 472802
rect 216588 472738 216640 472744
rect 215852 464364 215904 464370
rect 215852 464306 215904 464312
rect 215760 461644 215812 461650
rect 215760 461586 215812 461592
rect 215668 447364 215720 447370
rect 215668 447306 215720 447312
rect 215772 443972 215800 461586
rect 215864 447302 215892 464306
rect 215944 453416 215996 453422
rect 215944 453358 215996 453364
rect 215852 447296 215904 447302
rect 215852 447238 215904 447244
rect 215956 443972 215984 453358
rect 216496 447364 216548 447370
rect 216496 447306 216548 447312
rect 216312 447296 216364 447302
rect 216312 447238 216364 447244
rect 216128 447228 216180 447234
rect 216128 447170 216180 447176
rect 216140 443972 216168 447170
rect 216324 443972 216352 447238
rect 216508 443972 216536 447306
rect 216588 446548 216640 446554
rect 216588 446490 216640 446496
rect 216600 445126 216628 446490
rect 216588 445120 216640 445126
rect 216588 445062 216640 445068
rect 216692 443972 216720 482258
rect 216784 445126 216812 486406
rect 216956 483676 217008 483682
rect 216956 483618 217008 483624
rect 216864 463004 216916 463010
rect 216864 462946 216916 462952
rect 216772 445120 216824 445126
rect 216772 445062 216824 445068
rect 216876 443972 216904 462946
rect 216968 447250 216996 483618
rect 217140 475380 217192 475386
rect 217140 475322 217192 475328
rect 217152 447370 217180 475322
rect 217324 469872 217376 469878
rect 217324 469814 217376 469820
rect 217336 460934 217364 469814
rect 217508 465792 217560 465798
rect 217508 465734 217560 465740
rect 217520 460934 217548 465734
rect 217336 460906 217456 460934
rect 217520 460906 218008 460934
rect 217324 451920 217376 451926
rect 217324 451862 217376 451868
rect 217140 447364 217192 447370
rect 217140 447306 217192 447312
rect 216968 447222 217272 447250
rect 217048 444644 217100 444650
rect 217048 444586 217100 444592
rect 217060 443972 217088 444586
rect 217244 443972 217272 447222
rect 217336 444650 217364 451862
rect 217324 444644 217376 444650
rect 217324 444586 217376 444592
rect 217428 443972 217456 460906
rect 217600 447364 217652 447370
rect 217600 447306 217652 447312
rect 217612 443972 217640 447306
rect 217784 445120 217836 445126
rect 217784 445062 217836 445068
rect 217796 443972 217824 445062
rect 217980 443972 218008 460906
rect 218072 447370 218100 489126
rect 220084 488096 220136 488102
rect 220084 488038 220136 488044
rect 219808 487960 219860 487966
rect 219808 487902 219860 487908
rect 218244 478168 218296 478174
rect 218244 478110 218296 478116
rect 218152 476876 218204 476882
rect 218152 476818 218204 476824
rect 218060 447364 218112 447370
rect 218060 447306 218112 447312
rect 218164 443972 218192 476818
rect 218256 447302 218284 478110
rect 219624 468648 219676 468654
rect 219624 468590 219676 468596
rect 218336 468580 218388 468586
rect 218336 468522 218388 468528
rect 218244 447296 218296 447302
rect 218244 447238 218296 447244
rect 218348 443972 218376 468522
rect 218428 467220 218480 467226
rect 218428 467162 218480 467168
rect 218440 460934 218468 467162
rect 218440 460906 218560 460934
rect 218532 443972 218560 460906
rect 218612 460352 218664 460358
rect 218612 460294 218664 460300
rect 218624 445126 218652 460294
rect 219072 454708 219124 454714
rect 219072 454650 219124 454656
rect 218796 447704 218848 447710
rect 218796 447646 218848 447652
rect 218808 447302 218836 447646
rect 218888 447364 218940 447370
rect 218888 447306 218940 447312
rect 218704 447296 218756 447302
rect 218704 447238 218756 447244
rect 218796 447296 218848 447302
rect 218796 447238 218848 447244
rect 218612 445120 218664 445126
rect 218612 445062 218664 445068
rect 218716 443972 218744 447238
rect 218900 443972 218928 447306
rect 219084 443972 219112 454650
rect 219164 447772 219216 447778
rect 219164 447714 219216 447720
rect 219176 447438 219204 447714
rect 219440 447704 219492 447710
rect 219440 447646 219492 447652
rect 219164 447432 219216 447438
rect 219164 447374 219216 447380
rect 219348 445800 219400 445806
rect 219348 445742 219400 445748
rect 219256 445120 219308 445126
rect 219256 445062 219308 445068
rect 219268 443972 219296 445062
rect 219360 445058 219388 445742
rect 219348 445052 219400 445058
rect 219348 444994 219400 445000
rect 219452 443972 219480 447646
rect 219636 443972 219664 468590
rect 219716 463208 219768 463214
rect 219716 463150 219768 463156
rect 219728 452334 219756 463150
rect 219716 452328 219768 452334
rect 219716 452270 219768 452276
rect 219820 445040 219848 487902
rect 219900 461848 219952 461854
rect 219900 461790 219952 461796
rect 219912 447710 219940 461790
rect 220096 460934 220124 488038
rect 230572 488028 230624 488034
rect 230572 487970 230624 487976
rect 228364 487484 228416 487490
rect 228364 487426 228416 487432
rect 226984 487416 227036 487422
rect 226984 487358 227036 487364
rect 222844 487280 222896 487286
rect 220726 487248 220782 487257
rect 222844 487222 222896 487228
rect 226246 487248 226302 487257
rect 220726 487183 220782 487192
rect 220740 476814 220768 487183
rect 221464 484424 221516 484430
rect 221464 484366 221516 484372
rect 220728 476808 220780 476814
rect 220728 476750 220780 476756
rect 221372 467288 221424 467294
rect 221372 467230 221424 467236
rect 220096 460906 220216 460934
rect 219992 452328 220044 452334
rect 219992 452270 220044 452276
rect 219900 447704 219952 447710
rect 219900 447646 219952 447652
rect 219820 445012 219940 445040
rect 219912 444374 219940 445012
rect 219820 444346 219940 444374
rect 219820 443972 219848 444346
rect 220004 443972 220032 452270
rect 220084 445392 220136 445398
rect 220084 445334 220136 445340
rect 220096 444718 220124 445334
rect 220084 444712 220136 444718
rect 220084 444654 220136 444660
rect 220188 443972 220216 460906
rect 221004 458856 221056 458862
rect 221004 458798 221056 458804
rect 220820 457564 220872 457570
rect 220820 457506 220872 457512
rect 220728 451988 220780 451994
rect 220728 451930 220780 451936
rect 220360 446480 220412 446486
rect 220360 446422 220412 446428
rect 220372 443972 220400 446422
rect 220544 446412 220596 446418
rect 220544 446354 220596 446360
rect 220556 443972 220584 446354
rect 220740 443972 220768 451930
rect 220832 445126 220860 457506
rect 221016 447574 221044 458798
rect 221384 451274 221412 467230
rect 221476 451314 221504 484366
rect 221556 461712 221608 461718
rect 221556 461654 221608 461660
rect 221108 451246 221412 451274
rect 221464 451308 221516 451314
rect 221464 451250 221516 451256
rect 221004 447568 221056 447574
rect 221004 447510 221056 447516
rect 221108 447250 221136 451246
rect 221568 447250 221596 461654
rect 222016 457496 222068 457502
rect 222016 457438 222068 457444
rect 221740 453484 221792 453490
rect 221740 453426 221792 453432
rect 221648 448248 221700 448254
rect 221648 448190 221700 448196
rect 220924 447222 221136 447250
rect 221476 447222 221596 447250
rect 220820 445120 220872 445126
rect 220820 445062 220872 445068
rect 220924 443972 220952 447222
rect 221096 445392 221148 445398
rect 221096 445334 221148 445340
rect 221108 443972 221136 445334
rect 221280 445120 221332 445126
rect 221280 445062 221332 445068
rect 221292 443972 221320 445062
rect 221476 443972 221504 447222
rect 221660 446758 221688 448190
rect 221648 446752 221700 446758
rect 221648 446694 221700 446700
rect 221660 443972 221688 446694
rect 221752 445398 221780 453426
rect 221832 447568 221884 447574
rect 221832 447510 221884 447516
rect 221740 445392 221792 445398
rect 221740 445334 221792 445340
rect 221844 443972 221872 447510
rect 222028 443972 222056 457438
rect 222752 448588 222804 448594
rect 222752 448530 222804 448536
rect 222200 448520 222252 448526
rect 222200 448462 222252 448468
rect 222212 443972 222240 448462
rect 222384 448044 222436 448050
rect 222384 447986 222436 447992
rect 222396 443972 222424 447986
rect 222568 447976 222620 447982
rect 222568 447918 222620 447924
rect 222580 443972 222608 447918
rect 222764 443972 222792 448530
rect 222856 448390 222884 487222
rect 226246 487183 226302 487192
rect 224316 472728 224368 472734
rect 224316 472670 224368 472676
rect 223764 468512 223816 468518
rect 223764 468454 223816 468460
rect 222936 457292 222988 457298
rect 222936 457234 222988 457240
rect 222948 448526 222976 457234
rect 223028 456952 223080 456958
rect 223028 456894 223080 456900
rect 223040 449886 223068 456894
rect 223776 451274 223804 468454
rect 224224 464432 224276 464438
rect 224224 464374 224276 464380
rect 224040 460284 224092 460290
rect 224040 460226 224092 460232
rect 223856 456816 223908 456822
rect 223856 456758 223908 456764
rect 223684 451246 223804 451274
rect 223028 449880 223080 449886
rect 223028 449822 223080 449828
rect 223040 448594 223068 449822
rect 223120 449200 223172 449206
rect 223120 449142 223172 449148
rect 223028 448588 223080 448594
rect 223028 448530 223080 448536
rect 222936 448520 222988 448526
rect 222936 448462 222988 448468
rect 222844 448384 222896 448390
rect 222844 448326 222896 448332
rect 222936 448180 222988 448186
rect 222936 448122 222988 448128
rect 222948 443972 222976 448122
rect 223132 443972 223160 449142
rect 223488 448112 223540 448118
rect 223488 448054 223540 448060
rect 223304 447908 223356 447914
rect 223304 447850 223356 447856
rect 223316 446593 223344 447850
rect 223302 446584 223358 446593
rect 223302 446519 223358 446528
rect 223316 443972 223344 446519
rect 223500 443972 223528 448054
rect 223684 443972 223712 451246
rect 223868 443972 223896 456758
rect 224052 443972 224080 460226
rect 224236 451274 224264 464374
rect 224328 456822 224356 472670
rect 224500 471300 224552 471306
rect 224500 471242 224552 471248
rect 224512 460934 224540 471242
rect 224684 469940 224736 469946
rect 224684 469882 224736 469888
rect 224512 460906 224632 460934
rect 224316 456816 224368 456822
rect 224316 456758 224368 456764
rect 224236 451246 224448 451274
rect 224420 448633 224448 451246
rect 224406 448624 224462 448633
rect 224406 448559 224462 448568
rect 224224 445120 224276 445126
rect 224224 445062 224276 445068
rect 224236 443972 224264 445062
rect 224420 443972 224448 448559
rect 224604 443972 224632 460906
rect 224696 445126 224724 469882
rect 225604 462392 225656 462398
rect 225604 462334 225656 462340
rect 224776 447840 224828 447846
rect 224776 447782 224828 447788
rect 224684 445120 224736 445126
rect 224684 445062 224736 445068
rect 224788 443972 224816 447782
rect 225616 446894 225644 462334
rect 225694 454064 225750 454073
rect 225694 453999 225750 454008
rect 224960 446888 225012 446894
rect 224960 446830 225012 446836
rect 225604 446888 225656 446894
rect 225604 446830 225656 446836
rect 224972 446010 225000 446830
rect 225512 446616 225564 446622
rect 225512 446558 225564 446564
rect 224960 446004 225012 446010
rect 224960 445946 225012 445952
rect 224972 443972 225000 445946
rect 225144 445800 225196 445806
rect 225144 445742 225196 445748
rect 225156 443972 225184 445742
rect 225524 444145 225552 446558
rect 225708 445262 225736 453999
rect 226260 447846 226288 487183
rect 226996 448254 227024 487358
rect 227352 457496 227404 457502
rect 227352 457438 227404 457444
rect 226984 448248 227036 448254
rect 226984 448190 227036 448196
rect 226248 447840 226300 447846
rect 226248 447782 226300 447788
rect 227168 446548 227220 446554
rect 227168 446490 227220 446496
rect 226064 446140 226116 446146
rect 226064 446082 226116 446088
rect 225696 445256 225748 445262
rect 225696 445198 225748 445204
rect 225510 444136 225566 444145
rect 225510 444071 225566 444080
rect 225524 443972 225552 444071
rect 225708 443972 225736 445198
rect 226076 443972 226104 446082
rect 226984 446072 227036 446078
rect 226984 446014 227036 446020
rect 226246 445904 226302 445913
rect 226246 445839 226302 445848
rect 226260 445194 226288 445839
rect 226800 445324 226852 445330
rect 226800 445266 226852 445272
rect 226248 445188 226300 445194
rect 226248 445130 226300 445136
rect 226260 443972 226288 445130
rect 226706 444136 226762 444145
rect 226706 444071 226762 444080
rect 226524 443896 226576 443902
rect 226524 443838 226576 443844
rect 220452 443760 220504 443766
rect 226536 443748 226564 443838
rect 220452 443702 220504 443708
rect 225248 443720 225368 443748
rect 220464 443630 220492 443702
rect 220452 443624 220504 443630
rect 220452 443566 220504 443572
rect 211066 443456 211122 443465
rect 200948 443420 201000 443426
rect 211066 443391 211122 443400
rect 212354 443456 212410 443465
rect 212354 443391 212410 443400
rect 213642 443456 213698 443465
rect 225248 443426 225276 443720
rect 225340 443700 225368 443720
rect 225800 443720 225920 443748
rect 226352 443737 226472 443748
rect 225800 443494 225828 443720
rect 225892 443700 225920 443720
rect 226338 443728 226472 443737
rect 226394 443720 226472 443728
rect 226536 443720 226656 443748
rect 226720 443737 226748 444071
rect 226812 443972 226840 445266
rect 226996 443972 227024 446014
rect 227180 443972 227208 446490
rect 227364 444922 227392 457438
rect 228376 451246 228404 487426
rect 229744 487348 229796 487354
rect 229744 487290 229796 487296
rect 228456 457224 228508 457230
rect 228456 457166 228508 457172
rect 228364 451240 228416 451246
rect 228364 451182 228416 451188
rect 227536 446820 227588 446826
rect 227536 446762 227588 446768
rect 227352 444916 227404 444922
rect 227352 444858 227404 444864
rect 227364 443972 227392 444858
rect 227548 443972 227576 446762
rect 227720 445868 227772 445874
rect 227720 445810 227772 445816
rect 227732 443972 227760 445810
rect 228468 445738 228496 457166
rect 228548 457088 228600 457094
rect 228548 457030 228600 457036
rect 227904 445732 227956 445738
rect 227904 445674 227956 445680
rect 228456 445732 228508 445738
rect 228456 445674 228508 445680
rect 227916 444582 227944 445674
rect 228560 445618 228588 457030
rect 229756 449818 229784 487290
rect 229836 476808 229888 476814
rect 229836 476750 229888 476756
rect 229744 449812 229796 449818
rect 229744 449754 229796 449760
rect 229742 446720 229798 446729
rect 228640 446684 228692 446690
rect 229742 446655 229798 446664
rect 228640 446626 228692 446632
rect 228468 445590 228588 445618
rect 228468 444854 228496 445590
rect 228456 444848 228508 444854
rect 228456 444790 228508 444796
rect 227904 444576 227956 444582
rect 227904 444518 227956 444524
rect 227916 443972 227944 444518
rect 228468 443972 228496 444790
rect 228652 443972 228680 446626
rect 229190 446448 229246 446457
rect 229190 446383 229246 446392
rect 228824 445936 228876 445942
rect 228824 445878 228876 445884
rect 228836 443972 228864 445878
rect 229008 444440 229060 444446
rect 229008 444382 229060 444388
rect 229020 443972 229048 444382
rect 229204 443972 229232 446383
rect 229374 446040 229430 446049
rect 229374 445975 229430 445984
rect 229388 443972 229416 445975
rect 229560 445324 229612 445330
rect 229560 445266 229612 445272
rect 229572 444088 229600 445266
rect 229480 444060 229600 444088
rect 229480 443766 229508 444060
rect 229572 443972 229600 444060
rect 229756 443972 229784 446655
rect 229848 445874 229876 476750
rect 229928 475448 229980 475454
rect 229928 475390 229980 475396
rect 229940 446418 229968 475390
rect 230584 460934 230612 487970
rect 232596 487892 232648 487898
rect 232596 487834 232648 487840
rect 232504 487824 232556 487830
rect 232504 487766 232556 487772
rect 231766 487248 231822 487257
rect 231766 487183 231822 487192
rect 231492 464500 231544 464506
rect 231492 464442 231544 464448
rect 230756 463072 230808 463078
rect 230756 463014 230808 463020
rect 230768 460934 230796 463014
rect 231504 460934 231532 464442
rect 230584 460906 230704 460934
rect 230768 460906 231256 460934
rect 231504 460906 231624 460934
rect 230676 451058 230704 460906
rect 230676 451030 231072 451058
rect 230848 450968 230900 450974
rect 230848 450910 230900 450916
rect 230112 449948 230164 449954
rect 230112 449890 230164 449896
rect 229928 446412 229980 446418
rect 229928 446354 229980 446360
rect 229836 445868 229888 445874
rect 229836 445810 229888 445816
rect 229848 444060 229968 444088
rect 229468 443760 229520 443766
rect 226444 443700 226472 443720
rect 226628 443700 226656 443720
rect 226706 443728 226762 443737
rect 226338 443663 226394 443672
rect 226706 443663 226762 443672
rect 228008 443720 228128 443748
rect 225788 443488 225840 443494
rect 225788 443430 225840 443436
rect 228008 443426 228036 443720
rect 228100 443700 228128 443720
rect 228192 443720 228312 443748
rect 228192 443562 228220 443720
rect 228284 443700 228312 443720
rect 229468 443702 229520 443708
rect 229848 443698 229876 444060
rect 229940 443972 229968 444060
rect 230124 443972 230152 449890
rect 230664 446412 230716 446418
rect 230664 446354 230716 446360
rect 230480 444576 230532 444582
rect 230480 444518 230532 444524
rect 230308 444060 230428 444088
rect 230308 443972 230336 444060
rect 229836 443692 229888 443698
rect 229836 443634 229888 443640
rect 228180 443556 228232 443562
rect 228180 443498 228232 443504
rect 230400 443426 230428 444060
rect 230492 443972 230520 444518
rect 230676 443972 230704 446354
rect 230860 443972 230888 450910
rect 231044 443972 231072 451030
rect 231228 443972 231256 460906
rect 231596 459474 231624 460906
rect 231584 459468 231636 459474
rect 231584 459410 231636 459416
rect 231400 446072 231452 446078
rect 231400 446014 231452 446020
rect 231412 443972 231440 446014
rect 231596 443972 231624 459410
rect 231674 448760 231730 448769
rect 231674 448695 231730 448704
rect 231688 446026 231716 448695
rect 231780 447914 231808 487183
rect 232042 454336 232098 454345
rect 232042 454271 232098 454280
rect 231952 448384 232004 448390
rect 231952 448326 232004 448332
rect 231768 447908 231820 447914
rect 231768 447850 231820 447856
rect 231688 445998 231808 446026
rect 231780 443972 231808 445998
rect 231964 443972 231992 448326
rect 232056 447098 232084 454271
rect 232134 454200 232190 454209
rect 232134 454135 232190 454144
rect 232044 447092 232096 447098
rect 232044 447034 232096 447040
rect 232148 443972 232176 454135
rect 232516 448390 232544 487766
rect 232608 449138 232636 487834
rect 235906 487248 235962 487257
rect 235906 487183 235962 487192
rect 241426 487248 241482 487257
rect 244646 487248 244702 487257
rect 241426 487183 241482 487192
rect 244280 487212 244332 487218
rect 235264 486532 235316 486538
rect 235264 486474 235316 486480
rect 234620 482384 234672 482390
rect 234620 482326 234672 482332
rect 234632 451994 234660 482326
rect 235276 477494 235304 486474
rect 235264 477488 235316 477494
rect 235264 477430 235316 477436
rect 235276 476134 235304 477430
rect 234804 476128 234856 476134
rect 234804 476070 234856 476076
rect 235264 476128 235316 476134
rect 235264 476070 235316 476076
rect 234816 460934 234844 476070
rect 235920 473074 235948 487183
rect 238024 486600 238076 486606
rect 238024 486542 238076 486548
rect 236092 482384 236144 482390
rect 236092 482326 236144 482332
rect 235908 473068 235960 473074
rect 235908 473010 235960 473016
rect 235540 472796 235592 472802
rect 235540 472738 235592 472744
rect 235552 460934 235580 472738
rect 236000 472728 236052 472734
rect 236000 472670 236052 472676
rect 234816 460906 234936 460934
rect 235552 460906 235856 460934
rect 234620 451988 234672 451994
rect 234620 451930 234672 451936
rect 233976 451308 234028 451314
rect 233976 451250 234028 451256
rect 233424 450832 233476 450838
rect 233424 450774 233476 450780
rect 232688 449744 232740 449750
rect 232688 449686 232740 449692
rect 232596 449132 232648 449138
rect 232596 449074 232648 449080
rect 232504 448384 232556 448390
rect 232504 448326 232556 448332
rect 232608 447930 232636 449074
rect 232700 448390 232728 449686
rect 233056 449064 233108 449070
rect 233056 449006 233108 449012
rect 233068 448458 233096 449006
rect 233056 448452 233108 448458
rect 233056 448394 233108 448400
rect 232688 448384 232740 448390
rect 232688 448326 232740 448332
rect 232332 447902 232636 447930
rect 232332 443972 232360 447902
rect 232504 447092 232556 447098
rect 232504 447034 232556 447040
rect 232516 443972 232544 447034
rect 232700 443972 232728 448326
rect 232872 445800 232924 445806
rect 232872 445742 232924 445748
rect 232884 443972 232912 445742
rect 233068 443972 233096 448394
rect 233436 448186 233464 450774
rect 233792 450764 233844 450770
rect 233792 450706 233844 450712
rect 233804 448322 233832 450706
rect 233792 448316 233844 448322
rect 233792 448258 233844 448264
rect 233424 448180 233476 448186
rect 233424 448122 233476 448128
rect 233240 446412 233292 446418
rect 233240 446354 233292 446360
rect 233252 443972 233280 446354
rect 233436 443972 233464 448122
rect 233804 443972 233832 448258
rect 233988 443972 234016 451250
rect 234252 450900 234304 450906
rect 234252 450842 234304 450848
rect 234068 450696 234120 450702
rect 234068 450638 234120 450644
rect 234080 449857 234108 450638
rect 234264 449886 234292 450842
rect 234252 449880 234304 449886
rect 234066 449848 234122 449857
rect 234122 449806 234200 449834
rect 234252 449822 234304 449828
rect 234528 449880 234580 449886
rect 234528 449822 234580 449828
rect 234066 449783 234122 449792
rect 234172 443972 234200 449806
rect 234344 446140 234396 446146
rect 234344 446082 234396 446088
rect 234356 443972 234384 446082
rect 234540 443972 234568 449822
rect 234712 445188 234764 445194
rect 234712 445130 234764 445136
rect 234724 443972 234752 445130
rect 234908 443972 234936 460906
rect 235080 456000 235132 456006
rect 235080 455942 235132 455948
rect 235092 443972 235120 455942
rect 235356 454844 235408 454850
rect 235356 454786 235408 454792
rect 235264 454776 235316 454782
rect 235264 454718 235316 454724
rect 235276 443972 235304 454718
rect 235368 445194 235396 454786
rect 235632 451988 235684 451994
rect 235632 451930 235684 451936
rect 235356 445188 235408 445194
rect 235356 445130 235408 445136
rect 235448 444848 235500 444854
rect 235448 444790 235500 444796
rect 235460 443972 235488 444790
rect 235644 443972 235672 451930
rect 235828 443972 235856 460906
rect 236012 443972 236040 472670
rect 236104 460934 236132 482326
rect 236552 475516 236604 475522
rect 236552 475458 236604 475464
rect 236276 475448 236328 475454
rect 236276 475390 236328 475396
rect 236104 460906 236224 460934
rect 236196 443972 236224 460906
rect 236288 445194 236316 475390
rect 236564 460902 236592 475458
rect 237748 474088 237800 474094
rect 237748 474030 237800 474036
rect 237564 473340 237616 473346
rect 237564 473282 237616 473288
rect 237472 471300 237524 471306
rect 237472 471242 237524 471248
rect 236552 460896 236604 460902
rect 236552 460838 236604 460844
rect 236368 457156 236420 457162
rect 236368 457098 236420 457104
rect 236276 445188 236328 445194
rect 236276 445130 236328 445136
rect 236380 443972 236408 457098
rect 236564 443972 236592 460838
rect 236920 449268 236972 449274
rect 236920 449210 236972 449216
rect 236736 447976 236788 447982
rect 236736 447918 236788 447924
rect 236748 443972 236776 447918
rect 236932 443972 236960 449210
rect 237104 445868 237156 445874
rect 237104 445810 237156 445816
rect 237116 443972 237144 445810
rect 237288 445188 237340 445194
rect 237288 445130 237340 445136
rect 237300 443972 237328 445130
rect 237484 443972 237512 471242
rect 237576 452606 237604 473282
rect 237760 460934 237788 474030
rect 238036 473346 238064 486542
rect 239404 485240 239456 485246
rect 239404 485182 239456 485188
rect 238852 479664 238904 479670
rect 238852 479606 238904 479612
rect 238024 473340 238076 473346
rect 238024 473282 238076 473288
rect 237760 460906 238616 460934
rect 237748 455592 237800 455598
rect 237748 455534 237800 455540
rect 237564 452600 237616 452606
rect 237564 452542 237616 452548
rect 237760 444374 237788 455534
rect 237840 452600 237892 452606
rect 237840 452542 237892 452548
rect 237668 444346 237788 444374
rect 237668 443972 237696 444346
rect 237852 443972 237880 452542
rect 238208 449336 238260 449342
rect 238208 449278 238260 449284
rect 238022 444136 238078 444145
rect 238022 444071 238078 444080
rect 238036 443972 238064 444071
rect 238220 443972 238248 449278
rect 238392 447840 238444 447846
rect 238392 447782 238444 447788
rect 238404 443972 238432 447782
rect 238588 443972 238616 460906
rect 238760 445188 238812 445194
rect 238760 445130 238812 445136
rect 238772 443972 238800 445130
rect 238864 445126 238892 479606
rect 239036 468512 239088 468518
rect 239036 468454 239088 468460
rect 239048 451994 239076 468454
rect 239220 464432 239272 464438
rect 239220 464374 239272 464380
rect 239128 459536 239180 459542
rect 239128 459478 239180 459484
rect 239036 451988 239088 451994
rect 239036 451930 239088 451936
rect 238944 446480 238996 446486
rect 238944 446422 238996 446428
rect 238852 445120 238904 445126
rect 238852 445062 238904 445068
rect 238956 443972 238984 446422
rect 239140 443972 239168 459478
rect 239232 445194 239260 464374
rect 239416 459542 239444 485182
rect 240876 479732 240928 479738
rect 240876 479674 240928 479680
rect 240784 479596 240836 479602
rect 240784 479538 240836 479544
rect 240324 469940 240376 469946
rect 240324 469882 240376 469888
rect 239496 467152 239548 467158
rect 239496 467094 239548 467100
rect 239404 459536 239456 459542
rect 239404 459478 239456 459484
rect 239404 448316 239456 448322
rect 239404 448258 239456 448264
rect 239416 448118 239444 448258
rect 239404 448112 239456 448118
rect 239404 448054 239456 448060
rect 239312 445936 239364 445942
rect 239312 445878 239364 445884
rect 239220 445188 239272 445194
rect 239220 445130 239272 445136
rect 239324 443972 239352 445878
rect 239508 443972 239536 467094
rect 240336 451994 240364 469882
rect 240508 463140 240560 463146
rect 240508 463082 240560 463088
rect 240048 451988 240100 451994
rect 240048 451930 240100 451936
rect 240324 451988 240376 451994
rect 240324 451930 240376 451936
rect 239680 447908 239732 447914
rect 239680 447850 239732 447856
rect 239692 443972 239720 447850
rect 239864 445120 239916 445126
rect 239864 445062 239916 445068
rect 239876 443972 239904 445062
rect 240060 443972 240088 451930
rect 240416 448384 240468 448390
rect 240416 448326 240468 448332
rect 240428 448254 240456 448326
rect 240416 448248 240468 448254
rect 240416 448190 240468 448196
rect 240232 444916 240284 444922
rect 240232 444858 240284 444864
rect 240244 443972 240272 444858
rect 240428 443972 240456 448190
rect 240520 445194 240548 463082
rect 240796 448390 240824 479538
rect 240784 448384 240836 448390
rect 240784 448326 240836 448332
rect 240600 447568 240652 447574
rect 240600 447510 240652 447516
rect 240508 445188 240560 445194
rect 240508 445130 240560 445136
rect 240612 443972 240640 447510
rect 240888 447134 240916 479674
rect 241440 478990 241468 487183
rect 244646 487183 244702 487192
rect 249798 487248 249854 487257
rect 249798 487183 249854 487192
rect 244280 487154 244332 487160
rect 243820 485852 243872 485858
rect 243820 485794 243872 485800
rect 242164 483744 242216 483750
rect 242164 483686 242216 483692
rect 241428 478984 241480 478990
rect 241428 478926 241480 478932
rect 242176 474706 242204 483686
rect 243544 481092 243596 481098
rect 243544 481034 243596 481040
rect 242256 478984 242308 478990
rect 242256 478926 242308 478932
rect 241612 474700 241664 474706
rect 241612 474642 241664 474648
rect 242164 474700 242216 474706
rect 242164 474642 242216 474648
rect 240968 473068 241020 473074
rect 240968 473010 241020 473016
rect 240796 447106 240916 447134
rect 240796 443972 240824 447106
rect 240980 443972 241008 473010
rect 241624 460934 241652 474642
rect 242072 461780 242124 461786
rect 242072 461722 242124 461728
rect 241796 461712 241848 461718
rect 241796 461654 241848 461660
rect 241624 460906 241744 460934
rect 241336 451988 241388 451994
rect 241336 451930 241388 451936
rect 241152 445188 241204 445194
rect 241152 445130 241204 445136
rect 241164 443972 241192 445130
rect 241348 443972 241376 451930
rect 241520 449200 241572 449206
rect 241520 449142 241572 449148
rect 241532 443972 241560 449142
rect 241716 443972 241744 460906
rect 241808 445194 241836 461654
rect 241888 447636 241940 447642
rect 241888 447578 241940 447584
rect 241796 445188 241848 445194
rect 241796 445130 241848 445136
rect 241900 443972 241928 447578
rect 242084 443972 242112 461722
rect 242268 443972 242296 478926
rect 243360 465860 243412 465866
rect 243360 465802 243412 465808
rect 243084 465724 243136 465730
rect 243084 465666 243136 465672
rect 242992 449812 243044 449818
rect 242992 449754 243044 449760
rect 242624 445868 242676 445874
rect 242624 445810 242676 445816
rect 242440 445188 242492 445194
rect 242440 445130 242492 445136
rect 242452 443972 242480 445130
rect 242636 443972 242664 445810
rect 243004 443972 243032 449754
rect 243096 445194 243124 465666
rect 243176 452396 243228 452402
rect 243176 452338 243228 452344
rect 243084 445188 243136 445194
rect 243084 445130 243136 445136
rect 243188 443972 243216 452338
rect 243372 443972 243400 465802
rect 243556 449818 243584 481034
rect 243636 476808 243688 476814
rect 243636 476750 243688 476756
rect 243544 449812 243596 449818
rect 243544 449754 243596 449760
rect 243648 449392 243676 476750
rect 243464 449364 243676 449392
rect 243464 445874 243492 449364
rect 243832 447134 243860 485794
rect 244292 484362 244320 487154
rect 244660 485858 244688 487183
rect 249812 486674 249840 487183
rect 246488 486668 246540 486674
rect 246488 486610 246540 486616
rect 249800 486668 249852 486674
rect 249800 486610 249852 486616
rect 244924 486600 244976 486606
rect 244924 486542 244976 486548
rect 244648 485852 244700 485858
rect 244648 485794 244700 485800
rect 244280 484356 244332 484362
rect 244280 484298 244332 484304
rect 244292 480254 244320 484298
rect 244292 480226 244412 480254
rect 244280 451240 244332 451246
rect 244280 451182 244332 451188
rect 244292 450702 244320 451182
rect 244280 450696 244332 450702
rect 244280 450638 244332 450644
rect 243556 447106 243860 447134
rect 243452 445868 243504 445874
rect 243452 445810 243504 445816
rect 243556 443972 243584 447106
rect 243728 446888 243780 446894
rect 243728 446830 243780 446836
rect 243636 446480 243688 446486
rect 243636 446422 243688 446428
rect 243648 445942 243676 446422
rect 243636 445936 243688 445942
rect 243636 445878 243688 445884
rect 243740 443972 243768 446830
rect 243912 445188 243964 445194
rect 243912 445130 243964 445136
rect 243924 443972 243952 445130
rect 244096 445120 244148 445126
rect 244096 445062 244148 445068
rect 244108 443972 244136 445062
rect 244292 443972 244320 450638
rect 244384 445194 244412 480226
rect 244556 467152 244608 467158
rect 244556 467094 244608 467100
rect 244568 460934 244596 467094
rect 244568 460906 244872 460934
rect 244464 455728 244516 455734
rect 244464 455670 244516 455676
rect 244372 445188 244424 445194
rect 244372 445130 244424 445136
rect 244476 443972 244504 455670
rect 244648 449404 244700 449410
rect 244648 449346 244700 449352
rect 244660 443972 244688 449346
rect 244844 447250 244872 460906
rect 244936 450702 244964 486542
rect 245660 474156 245712 474162
rect 245660 474098 245712 474104
rect 245672 460934 245700 474098
rect 245672 460906 245792 460934
rect 244924 450696 244976 450702
rect 244924 450638 244976 450644
rect 245660 447840 245712 447846
rect 245660 447782 245712 447788
rect 244844 447222 245240 447250
rect 244832 446480 244884 446486
rect 244832 446422 244884 446428
rect 244844 445942 244872 446422
rect 244832 445936 244884 445942
rect 244832 445878 244884 445884
rect 245016 445868 245068 445874
rect 245016 445810 245068 445816
rect 244832 445800 244884 445806
rect 244832 445742 244884 445748
rect 244844 443972 244872 445742
rect 245028 443972 245056 445810
rect 245212 443972 245240 447222
rect 245672 447134 245700 447782
rect 245764 447250 245792 460906
rect 245844 460284 245896 460290
rect 245844 460226 245896 460232
rect 245856 447778 245884 460226
rect 246304 458380 246356 458386
rect 246304 458322 246356 458328
rect 246028 452056 246080 452062
rect 246028 451998 246080 452004
rect 245844 447772 245896 447778
rect 245844 447714 245896 447720
rect 246040 447710 246068 451998
rect 246120 449608 246172 449614
rect 246120 449550 246172 449556
rect 246028 447704 246080 447710
rect 246028 447646 246080 447652
rect 245764 447222 245976 447250
rect 245672 447106 245792 447134
rect 245660 445732 245712 445738
rect 245660 445674 245712 445680
rect 245568 445188 245620 445194
rect 245568 445130 245620 445136
rect 245474 444000 245530 444009
rect 245580 443972 245608 445130
rect 245474 443935 245530 443944
rect 245488 443884 245516 443935
rect 245396 443856 245516 443884
rect 245396 443836 245424 443856
rect 245672 443698 245700 445674
rect 245764 443972 245792 447106
rect 245948 443972 245976 447222
rect 246132 443972 246160 449550
rect 246316 447642 246344 458322
rect 246396 447772 246448 447778
rect 246396 447714 246448 447720
rect 246304 447636 246356 447642
rect 246304 447578 246356 447584
rect 246408 447250 246436 447714
rect 246500 447658 246528 486610
rect 248420 486532 248472 486538
rect 248420 486474 248472 486480
rect 247868 481024 247920 481030
rect 247868 480966 247920 480972
rect 246580 478236 246632 478242
rect 246580 478178 246632 478184
rect 246592 460934 246620 478178
rect 247880 460934 247908 480966
rect 246592 460906 246712 460934
rect 247880 460906 248092 460934
rect 246500 447630 246620 447658
rect 246408 447222 246528 447250
rect 246304 446616 246356 446622
rect 246304 446558 246356 446564
rect 246316 443972 246344 446558
rect 246500 443972 246528 447222
rect 246592 445806 246620 447630
rect 246684 446894 246712 460906
rect 247040 458856 247092 458862
rect 247040 458798 247092 458804
rect 247052 452402 247080 458798
rect 247132 457020 247184 457026
rect 247132 456962 247184 456968
rect 247040 452396 247092 452402
rect 247040 452338 247092 452344
rect 246764 449268 246816 449274
rect 246764 449210 246816 449216
rect 246672 446888 246724 446894
rect 246672 446830 246724 446836
rect 246580 445800 246632 445806
rect 246580 445742 246632 445748
rect 246776 445210 246804 449210
rect 247040 448588 247092 448594
rect 247040 448530 247092 448536
rect 246856 447704 246908 447710
rect 246856 447646 246908 447652
rect 246684 445182 246804 445210
rect 246684 443972 246712 445182
rect 246868 443972 246896 447646
rect 247052 443972 247080 448530
rect 247144 445398 247172 456962
rect 247316 452124 247368 452130
rect 247316 452066 247368 452072
rect 247224 449540 247276 449546
rect 247224 449482 247276 449488
rect 247132 445392 247184 445398
rect 247132 445334 247184 445340
rect 247236 443972 247264 449482
rect 247328 445194 247356 452066
rect 247776 451988 247828 451994
rect 247776 451930 247828 451936
rect 247408 449676 247460 449682
rect 247408 449618 247460 449624
rect 247316 445188 247368 445194
rect 247316 445130 247368 445136
rect 247420 443972 247448 449618
rect 247788 447250 247816 451930
rect 247788 447222 248000 447250
rect 247776 446888 247828 446894
rect 247776 446830 247828 446836
rect 247592 446548 247644 446554
rect 247592 446490 247644 446496
rect 247604 443972 247632 446490
rect 247788 443972 247816 446830
rect 247972 443972 248000 447222
rect 248064 445874 248092 460906
rect 248052 445868 248104 445874
rect 248052 445810 248104 445816
rect 248328 445392 248380 445398
rect 248328 445334 248380 445340
rect 248144 445188 248196 445194
rect 248144 445130 248196 445136
rect 248156 443972 248184 445130
rect 248340 443972 248368 445334
rect 248432 445194 248460 486474
rect 251180 483744 251232 483750
rect 251180 483686 251232 483692
rect 250812 481160 250864 481166
rect 250812 481102 250864 481108
rect 248512 478304 248564 478310
rect 248512 478246 248564 478252
rect 248420 445188 248472 445194
rect 248420 445130 248472 445136
rect 248524 443972 248552 478246
rect 250824 460934 250852 481102
rect 251192 460934 251220 483686
rect 250824 460906 251128 460934
rect 251192 460906 251680 460934
rect 249800 458924 249852 458930
rect 249800 458866 249852 458872
rect 249248 454912 249300 454918
rect 249248 454854 249300 454860
rect 248696 449404 248748 449410
rect 248696 449346 248748 449352
rect 248604 446752 248656 446758
rect 248604 446694 248656 446700
rect 248616 445058 248644 446694
rect 248604 445052 248656 445058
rect 248604 444994 248656 445000
rect 248708 443972 248736 449346
rect 248880 447908 248932 447914
rect 248880 447850 248932 447856
rect 248892 443972 248920 447850
rect 249064 445188 249116 445194
rect 249064 445130 249116 445136
rect 249076 443972 249104 445130
rect 249260 443972 249288 454854
rect 249432 449336 249484 449342
rect 249432 449278 249484 449284
rect 249444 443972 249472 449278
rect 249812 443972 249840 458866
rect 250536 455796 250588 455802
rect 250536 455738 250588 455744
rect 249984 449608 250036 449614
rect 249984 449550 250036 449556
rect 249892 445936 249944 445942
rect 249892 445878 249944 445884
rect 249628 443856 249748 443884
rect 249628 443836 249656 443856
rect 245660 443692 245712 443698
rect 245660 443634 245712 443640
rect 249720 443426 249748 443856
rect 249904 443766 249932 445878
rect 249996 443972 250024 449550
rect 250352 446956 250404 446962
rect 250352 446898 250404 446904
rect 250168 446820 250220 446826
rect 250168 446762 250220 446768
rect 250180 443972 250208 446762
rect 250364 443972 250392 446898
rect 250548 443972 250576 455738
rect 250720 449540 250772 449546
rect 250720 449482 250772 449488
rect 250732 443972 250760 449482
rect 250994 444000 251050 444009
rect 251100 443972 251128 460906
rect 251272 449676 251324 449682
rect 251272 449618 251324 449624
rect 251284 443972 251312 449618
rect 251456 446752 251508 446758
rect 251456 446694 251508 446700
rect 251468 443972 251496 446694
rect 251652 443972 251680 460906
rect 251824 458924 251876 458930
rect 251824 458866 251876 458872
rect 251836 447982 251864 458866
rect 252744 455932 252796 455938
rect 252744 455874 252796 455880
rect 251916 455864 251968 455870
rect 251916 455806 251968 455812
rect 251824 447976 251876 447982
rect 251824 447918 251876 447924
rect 251928 446418 251956 455806
rect 252560 449744 252612 449750
rect 252560 449686 252612 449692
rect 252008 449472 252060 449478
rect 252008 449414 252060 449420
rect 251916 446412 251968 446418
rect 251916 446354 251968 446360
rect 251824 445188 251876 445194
rect 251824 445130 251876 445136
rect 251836 443972 251864 445130
rect 252020 443972 252048 449414
rect 252376 448996 252428 449002
rect 252376 448938 252428 448944
rect 252192 448656 252244 448662
rect 252192 448598 252244 448604
rect 252204 443972 252232 448598
rect 252388 443972 252416 448938
rect 252572 443972 252600 449686
rect 252756 447250 252784 455874
rect 253296 452192 253348 452198
rect 253296 452134 253348 452140
rect 252756 447222 253152 447250
rect 252928 447092 252980 447098
rect 252928 447034 252980 447040
rect 252744 446684 252796 446690
rect 252744 446626 252796 446632
rect 252652 446480 252704 446486
rect 252652 446422 252704 446428
rect 250994 443935 251050 443944
rect 251008 443884 251036 443935
rect 250916 443856 251036 443884
rect 250916 443836 250944 443856
rect 252664 443834 252692 446422
rect 252756 443972 252784 446626
rect 252940 443972 252968 447034
rect 253124 443972 253152 447222
rect 253308 443972 253336 452134
rect 253478 444272 253534 444281
rect 253478 444207 253534 444216
rect 253492 443972 253520 444207
rect 253676 443972 253704 489194
rect 254952 485172 255004 485178
rect 254952 485114 255004 485120
rect 253940 485104 253992 485110
rect 253940 485046 253992 485052
rect 253952 460934 253980 485046
rect 253952 460906 254072 460934
rect 253848 449812 253900 449818
rect 253848 449754 253900 449760
rect 253860 443972 253888 449754
rect 254044 447250 254072 460906
rect 254584 452260 254636 452266
rect 254584 452202 254636 452208
rect 254044 447222 254256 447250
rect 254032 446412 254084 446418
rect 254032 446354 254084 446360
rect 254044 443972 254072 446354
rect 254228 443972 254256 447222
rect 254308 446004 254360 446010
rect 254308 445946 254360 445952
rect 254320 443902 254348 445946
rect 254398 444408 254454 444417
rect 254398 444343 254454 444352
rect 254412 443972 254440 444343
rect 254596 443972 254624 452202
rect 254768 450764 254820 450770
rect 254768 450706 254820 450712
rect 254780 443972 254808 450706
rect 254964 443972 254992 485114
rect 255872 452328 255924 452334
rect 255872 452270 255924 452276
rect 255688 450696 255740 450702
rect 255688 450638 255740 450644
rect 255412 450628 255464 450634
rect 255412 450570 255464 450576
rect 255320 450560 255372 450566
rect 255320 450502 255372 450508
rect 255136 449132 255188 449138
rect 255136 449074 255188 449080
rect 255148 443972 255176 449074
rect 255332 448254 255360 450502
rect 255424 449721 255452 450570
rect 255410 449712 255466 449721
rect 255410 449647 255466 449656
rect 255320 448248 255372 448254
rect 255320 448190 255372 448196
rect 255320 447024 255372 447030
rect 255320 446966 255372 446972
rect 255332 443972 255360 446966
rect 255502 446448 255558 446457
rect 255502 446383 255558 446392
rect 255412 446072 255464 446078
rect 255412 446014 255464 446020
rect 255424 444038 255452 446014
rect 255412 444032 255464 444038
rect 255412 443974 255464 443980
rect 255516 443972 255544 446383
rect 255596 446140 255648 446146
rect 255596 446082 255648 446088
rect 255608 443970 255636 446082
rect 255700 443972 255728 450638
rect 255884 443972 255912 452270
rect 256056 450832 256108 450838
rect 256056 450774 256108 450780
rect 256068 443972 256096 450774
rect 256422 449712 256478 449721
rect 256422 449647 256478 449656
rect 256240 448248 256292 448254
rect 256240 448190 256292 448196
rect 256252 443972 256280 448190
rect 256436 444145 256464 449647
rect 281000 447914 281028 597314
rect 281080 596760 281132 596766
rect 281080 596702 281132 596708
rect 281092 596222 281120 596702
rect 281540 596488 281592 596494
rect 281540 596430 281592 596436
rect 281552 596358 281580 596430
rect 281540 596352 281592 596358
rect 281540 596294 281592 596300
rect 281080 596216 281132 596222
rect 281080 596158 281132 596164
rect 281092 452062 281120 596158
rect 281552 452130 281580 596294
rect 282184 592680 282236 592686
rect 282184 592622 282236 592628
rect 281632 581664 281684 581670
rect 281632 581606 281684 581612
rect 281540 452124 281592 452130
rect 281540 452066 281592 452072
rect 281080 452056 281132 452062
rect 281080 451998 281132 452004
rect 281644 449410 281672 581606
rect 281724 580576 281776 580582
rect 281724 580518 281776 580524
rect 281632 449404 281684 449410
rect 281632 449346 281684 449352
rect 281736 449138 281764 580518
rect 281816 580508 281868 580514
rect 281816 580450 281868 580456
rect 281828 449818 281856 580450
rect 282092 580440 282144 580446
rect 282092 580382 282144 580388
rect 281908 580372 281960 580378
rect 281908 580314 281960 580320
rect 281816 449812 281868 449818
rect 281816 449754 281868 449760
rect 281920 449682 281948 580314
rect 282000 580304 282052 580310
rect 282000 580246 282052 580252
rect 281908 449676 281960 449682
rect 281908 449618 281960 449624
rect 282012 449614 282040 580246
rect 282104 449750 282132 580382
rect 282092 449744 282144 449750
rect 282092 449686 282144 449692
rect 282000 449608 282052 449614
rect 282000 449550 282052 449556
rect 281724 449132 281776 449138
rect 281724 449074 281776 449080
rect 280988 447908 281040 447914
rect 280988 447850 281040 447856
rect 282196 446894 282224 592622
rect 282276 587172 282328 587178
rect 282276 587114 282328 587120
rect 282288 446962 282316 587114
rect 282368 580304 282420 580310
rect 282368 580246 282420 580252
rect 282380 447098 282408 580246
rect 282932 463214 282960 702406
rect 300136 700534 300164 703520
rect 296076 700528 296128 700534
rect 296076 700470 296128 700476
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 293224 700460 293276 700466
rect 293224 700402 293276 700408
rect 291844 700392 291896 700398
rect 291844 700334 291896 700340
rect 283012 700324 283064 700330
rect 283012 700266 283064 700272
rect 283024 487966 283052 700266
rect 286324 696992 286376 696998
rect 286324 696934 286376 696940
rect 284576 597032 284628 597038
rect 284576 596974 284628 596980
rect 284392 596964 284444 596970
rect 284392 596906 284444 596912
rect 283196 596828 283248 596834
rect 283196 596770 283248 596776
rect 283104 596692 283156 596698
rect 283104 596634 283156 596640
rect 283116 596290 283144 596634
rect 283208 596630 283236 596770
rect 283196 596624 283248 596630
rect 283196 596566 283248 596572
rect 283104 596284 283156 596290
rect 283104 596226 283156 596232
rect 283012 487960 283064 487966
rect 283012 487902 283064 487908
rect 282920 463208 282972 463214
rect 282920 463150 282972 463156
rect 283116 449342 283144 596226
rect 283208 449546 283236 596566
rect 284300 596556 284352 596562
rect 284300 596498 284352 596504
rect 284312 596426 284340 596498
rect 284300 596420 284352 596426
rect 284300 596362 284352 596368
rect 283196 449540 283248 449546
rect 283196 449482 283248 449488
rect 284312 449478 284340 596362
rect 284404 596290 284432 596906
rect 284484 596896 284536 596902
rect 284484 596838 284536 596844
rect 284496 596358 284524 596838
rect 284588 596426 284616 596974
rect 284576 596420 284628 596426
rect 284576 596362 284628 596368
rect 284484 596352 284536 596358
rect 284484 596294 284536 596300
rect 284392 596284 284444 596290
rect 284392 596226 284444 596232
rect 284404 452334 284432 596226
rect 284392 452328 284444 452334
rect 284392 452270 284444 452276
rect 284496 452266 284524 596294
rect 284484 452260 284536 452266
rect 284484 452202 284536 452208
rect 284588 452198 284616 596362
rect 285036 590708 285088 590714
rect 285036 590650 285088 590656
rect 284944 588600 284996 588606
rect 284944 588542 284996 588548
rect 284576 452192 284628 452198
rect 284576 452134 284628 452140
rect 284300 449472 284352 449478
rect 284300 449414 284352 449420
rect 283104 449336 283156 449342
rect 283104 449278 283156 449284
rect 282368 447092 282420 447098
rect 282368 447034 282420 447040
rect 282276 446956 282328 446962
rect 282276 446898 282328 446904
rect 282184 446888 282236 446894
rect 282184 446830 282236 446836
rect 284956 446826 284984 588542
rect 285048 453422 285076 590650
rect 285036 453416 285088 453422
rect 285036 453358 285088 453364
rect 286336 451926 286364 696934
rect 289084 589960 289136 589966
rect 289084 589902 289136 589908
rect 287704 587240 287756 587246
rect 287704 587182 287756 587188
rect 286416 585880 286468 585886
rect 286416 585822 286468 585828
rect 286324 451920 286376 451926
rect 286324 451862 286376 451868
rect 286428 447030 286456 585822
rect 286416 447024 286468 447030
rect 286416 446966 286468 446972
rect 284944 446820 284996 446826
rect 284944 446762 284996 446768
rect 287716 446622 287744 587182
rect 287796 498840 287848 498846
rect 287796 498782 287848 498788
rect 287808 488034 287836 498782
rect 287796 488028 287848 488034
rect 287796 487970 287848 487976
rect 287704 446616 287756 446622
rect 287704 446558 287756 446564
rect 289096 446554 289124 589902
rect 289176 581664 289228 581670
rect 289176 581606 289228 581612
rect 289188 446758 289216 581606
rect 291856 461854 291884 700334
rect 291936 583024 291988 583030
rect 291936 582966 291988 582972
rect 291844 461848 291896 461854
rect 291844 461790 291896 461796
rect 289176 446752 289228 446758
rect 289176 446694 289228 446700
rect 291948 446690 291976 582966
rect 292028 488436 292080 488442
rect 292028 488378 292080 488384
rect 292040 449721 292068 488378
rect 293236 460358 293264 700402
rect 295984 700324 296036 700330
rect 295984 700266 296036 700272
rect 293868 526788 293920 526794
rect 293868 526730 293920 526736
rect 293880 488481 293908 526730
rect 293314 488472 293370 488481
rect 293314 488407 293370 488416
rect 293866 488472 293922 488481
rect 293866 488407 293922 488416
rect 293328 477494 293356 488407
rect 293880 488073 293908 488407
rect 293866 488064 293922 488073
rect 293866 487999 293922 488008
rect 293316 477488 293368 477494
rect 293316 477430 293368 477436
rect 293224 460352 293276 460358
rect 293224 460294 293276 460300
rect 293316 458312 293368 458318
rect 293316 458254 293368 458260
rect 293328 450838 293356 458254
rect 295996 454714 296024 700266
rect 296088 468654 296116 700470
rect 332520 700466 332548 703520
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364996 700330 365024 703520
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 397472 699718 397500 703520
rect 413664 700602 413692 703520
rect 405004 700596 405056 700602
rect 405004 700538 405056 700544
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 403624 700460 403676 700466
rect 403624 700402 403676 700408
rect 399484 700392 399536 700398
rect 399484 700334 399536 700340
rect 395344 699712 395396 699718
rect 395344 699654 395396 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 298006 636984 298062 636993
rect 298006 636919 298062 636928
rect 297178 635896 297234 635905
rect 297178 635831 297234 635840
rect 297086 610192 297142 610201
rect 297086 610127 297142 610136
rect 296994 608696 297050 608705
rect 296994 608631 297050 608640
rect 296902 517576 296958 517585
rect 296902 517511 296958 517520
rect 296916 488345 296944 517511
rect 297008 498846 297036 608631
rect 297100 500313 297128 610127
rect 297192 585818 297220 635831
rect 297914 634264 297970 634273
rect 297914 634199 297970 634208
rect 297730 633176 297786 633185
rect 297730 633111 297786 633120
rect 297454 631544 297510 631553
rect 297454 631479 297510 631488
rect 297364 600160 297416 600166
rect 297364 600102 297416 600108
rect 297272 598596 297324 598602
rect 297272 598538 297324 598544
rect 297180 585812 297232 585818
rect 297180 585754 297232 585760
rect 297192 526017 297220 585754
rect 297284 526794 297312 598538
rect 297272 526788 297324 526794
rect 297272 526730 297324 526736
rect 297178 526008 297234 526017
rect 297178 525943 297234 525952
rect 297086 500304 297142 500313
rect 297086 500239 297142 500248
rect 296996 498840 297048 498846
rect 296996 498782 297048 498788
rect 297100 488510 297128 500239
rect 297088 488504 297140 488510
rect 297088 488446 297140 488452
rect 296902 488336 296958 488345
rect 296902 488271 296958 488280
rect 296076 468648 296128 468654
rect 296076 468590 296128 468596
rect 296076 458652 296128 458658
rect 296076 458594 296128 458600
rect 295984 454708 296036 454714
rect 295984 454650 296036 454656
rect 293316 450832 293368 450838
rect 293316 450774 293368 450780
rect 293224 449948 293276 449954
rect 293224 449890 293276 449896
rect 292026 449712 292082 449721
rect 292026 449647 292082 449656
rect 291936 446684 291988 446690
rect 291936 446626 291988 446632
rect 289084 446548 289136 446554
rect 289084 446490 289136 446496
rect 256608 446480 256660 446486
rect 256608 446422 256660 446428
rect 256422 444136 256478 444145
rect 256422 444071 256478 444080
rect 256436 443972 256464 444071
rect 256620 443972 256648 446422
rect 256790 445768 256846 445777
rect 256790 445703 256846 445712
rect 256804 443972 256832 445703
rect 267004 445324 267056 445330
rect 267004 445266 267056 445272
rect 265900 445256 265952 445262
rect 265900 445198 265952 445204
rect 265716 444984 265768 444990
rect 265716 444926 265768 444932
rect 265622 444680 265678 444689
rect 265622 444615 265678 444624
rect 255596 443964 255648 443970
rect 255596 443906 255648 443912
rect 254308 443896 254360 443902
rect 254308 443838 254360 443844
rect 252652 443828 252704 443834
rect 252652 443770 252704 443776
rect 249892 443760 249944 443766
rect 249892 443702 249944 443708
rect 213642 443391 213698 443400
rect 225236 443420 225288 443426
rect 200948 443362 201000 443368
rect 225236 443362 225288 443368
rect 227996 443420 228048 443426
rect 227996 443362 228048 443368
rect 230388 443420 230440 443426
rect 233700 443420 233752 443426
rect 230388 443362 230440 443368
rect 233620 443380 233700 443408
rect 200960 306338 200988 443362
rect 233620 443292 233648 443380
rect 242900 443420 242952 443426
rect 233700 443362 233752 443368
rect 242820 443380 242900 443408
rect 242820 443292 242848 443380
rect 242900 443362 242952 443368
rect 249708 443420 249760 443426
rect 249708 443362 249760 443368
rect 205640 399152 205692 399158
rect 205640 399094 205692 399100
rect 210240 399152 210292 399158
rect 210240 399094 210292 399100
rect 203430 398848 203486 398857
rect 203430 398783 203486 398792
rect 202142 398440 202198 398449
rect 202142 398375 202198 398384
rect 201500 397316 201552 397322
rect 201500 397258 201552 397264
rect 200948 306332 201000 306338
rect 200948 306274 201000 306280
rect 200856 71732 200908 71738
rect 200856 71674 200908 71680
rect 200764 20664 200816 20670
rect 200764 20606 200816 20612
rect 200304 6656 200356 6662
rect 200304 6598 200356 6604
rect 200316 480 200344 6598
rect 201512 3398 201540 397258
rect 202156 181490 202184 398375
rect 203444 397497 203472 398783
rect 203706 398712 203762 398721
rect 203706 398647 203762 398656
rect 203522 398576 203578 398585
rect 203522 398511 203578 398520
rect 203430 397488 203486 397497
rect 203430 397423 203486 397432
rect 202880 394324 202932 394330
rect 202880 394266 202932 394272
rect 202144 181484 202196 181490
rect 202144 181426 202196 181432
rect 202892 16574 202920 394266
rect 202892 16546 203472 16574
rect 201592 5432 201644 5438
rect 201592 5374 201644 5380
rect 201500 3392 201552 3398
rect 201500 3334 201552 3340
rect 201604 2802 201632 5374
rect 202696 3392 202748 3398
rect 202696 3334 202748 3340
rect 201512 2774 201632 2802
rect 201512 480 201540 2774
rect 202708 480 202736 3334
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203536 4826 203564 398511
rect 203720 169046 203748 398647
rect 203708 169040 203760 169046
rect 203708 168982 203760 168988
rect 205652 16574 205680 399094
rect 207664 399084 207716 399090
rect 207664 399026 207716 399032
rect 206284 398812 206336 398818
rect 206284 398754 206336 398760
rect 205822 398712 205878 398721
rect 205822 398647 205878 398656
rect 205836 398449 205864 398647
rect 205822 398440 205878 398449
rect 205822 398375 205878 398384
rect 206296 86290 206324 398754
rect 207020 398404 207072 398410
rect 207020 398346 207072 398352
rect 206284 86284 206336 86290
rect 206284 86226 206336 86232
rect 205652 16546 206232 16574
rect 203524 4820 203576 4826
rect 203524 4762 203576 4768
rect 205088 4820 205140 4826
rect 205088 4762 205140 4768
rect 205100 480 205128 4762
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 398346
rect 207676 3670 207704 399026
rect 209872 398948 209924 398954
rect 209872 398890 209924 398896
rect 209884 398834 209912 398890
rect 210252 398886 210280 399094
rect 209792 398806 209912 398834
rect 210240 398880 210292 398886
rect 210240 398822 210292 398828
rect 207756 398676 207808 398682
rect 207756 398618 207808 398624
rect 207768 3806 207796 398618
rect 208400 398540 208452 398546
rect 208400 398482 208452 398488
rect 208032 398472 208084 398478
rect 208032 398414 208084 398420
rect 207848 397928 207900 397934
rect 207848 397870 207900 397876
rect 207860 83502 207888 397870
rect 207940 397860 207992 397866
rect 207940 397802 207992 397808
rect 207952 180130 207980 397802
rect 208044 340202 208072 398414
rect 208032 340196 208084 340202
rect 208032 340138 208084 340144
rect 207940 180124 207992 180130
rect 207940 180066 207992 180072
rect 207848 83496 207900 83502
rect 207848 83438 207900 83444
rect 208412 16574 208440 398482
rect 209320 398064 209372 398070
rect 209320 398006 209372 398012
rect 209136 397724 209188 397730
rect 209136 397666 209188 397672
rect 209044 397248 209096 397254
rect 209044 397190 209096 397196
rect 208412 16546 208624 16574
rect 207756 3800 207808 3806
rect 207756 3742 207808 3748
rect 207664 3664 207716 3670
rect 207664 3606 207716 3612
rect 208596 480 208624 16546
rect 209056 3874 209084 397190
rect 209148 333266 209176 397666
rect 209228 397656 209280 397662
rect 209228 397598 209280 397604
rect 209240 338774 209268 397598
rect 209332 363662 209360 398006
rect 209320 363656 209372 363662
rect 209320 363598 209372 363604
rect 209228 338768 209280 338774
rect 209228 338710 209280 338716
rect 209136 333260 209188 333266
rect 209136 333202 209188 333208
rect 209792 9674 209820 398806
rect 210344 397633 210372 400044
rect 210330 397624 210386 397633
rect 210330 397559 210386 397568
rect 210436 397497 210464 400044
rect 210422 397488 210478 397497
rect 210422 397423 210478 397432
rect 210422 397352 210478 397361
rect 210422 397287 210478 397296
rect 209870 396400 209926 396409
rect 209870 396335 209926 396344
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 396335
rect 210436 396074 210464 397287
rect 210344 396046 210464 396074
rect 210148 393916 210200 393922
rect 210148 393858 210200 393864
rect 209964 393848 210016 393854
rect 209964 393790 210016 393796
rect 209976 8974 210004 393790
rect 210056 392216 210108 392222
rect 210056 392158 210108 392164
rect 210068 9042 210096 392158
rect 210160 13122 210188 393858
rect 210344 391270 210372 396046
rect 210528 393854 210556 400044
rect 210620 393922 210648 400044
rect 210712 393990 210740 400044
rect 210700 393984 210752 393990
rect 210700 393926 210752 393932
rect 210608 393916 210660 393922
rect 210608 393858 210660 393864
rect 210516 393848 210568 393854
rect 210516 393790 210568 393796
rect 210804 391354 210832 400044
rect 210896 392222 210924 400044
rect 210884 392216 210936 392222
rect 210884 392158 210936 392164
rect 210436 391326 210832 391354
rect 210332 391264 210384 391270
rect 210332 391206 210384 391212
rect 210240 390584 210292 390590
rect 210240 390526 210292 390532
rect 210252 13190 210280 390526
rect 210332 390516 210384 390522
rect 210332 390458 210384 390464
rect 210344 177342 210372 390458
rect 210436 352578 210464 391326
rect 210516 391264 210568 391270
rect 210516 391206 210568 391212
rect 210424 352572 210476 352578
rect 210424 352514 210476 352520
rect 210528 351218 210556 391206
rect 210988 390590 211016 400044
rect 210976 390584 211028 390590
rect 210976 390526 211028 390532
rect 211080 390522 211108 400044
rect 211172 398313 211200 400044
rect 211158 398304 211214 398313
rect 211158 398239 211214 398248
rect 211158 397896 211214 397905
rect 211158 397831 211214 397840
rect 211172 396846 211200 397831
rect 211264 397769 211292 400044
rect 211250 397760 211306 397769
rect 211250 397695 211306 397704
rect 211356 397497 211384 400044
rect 211448 398313 211476 400044
rect 211434 398304 211490 398313
rect 211434 398239 211490 398248
rect 211436 398132 211488 398138
rect 211436 398074 211488 398080
rect 211342 397488 211398 397497
rect 211342 397423 211398 397432
rect 211160 396840 211212 396846
rect 211160 396782 211212 396788
rect 211448 395350 211476 398074
rect 211540 398041 211568 400044
rect 211526 398032 211582 398041
rect 211526 397967 211582 397976
rect 211632 397633 211660 400044
rect 211618 397624 211674 397633
rect 211618 397559 211674 397568
rect 211436 395344 211488 395350
rect 211436 395286 211488 395292
rect 211724 394040 211752 400044
rect 211816 398585 211844 400044
rect 211908 398721 211936 400044
rect 211894 398712 211950 398721
rect 211894 398647 211950 398656
rect 211896 398608 211948 398614
rect 211802 398576 211858 398585
rect 211896 398550 211948 398556
rect 211802 398511 211858 398520
rect 211802 397624 211858 397633
rect 211802 397559 211858 397568
rect 211356 394012 211752 394040
rect 211068 390516 211120 390522
rect 211068 390458 211120 390464
rect 210516 351212 210568 351218
rect 210516 351154 210568 351160
rect 210332 177336 210384 177342
rect 210332 177278 210384 177284
rect 211356 14482 211384 394012
rect 211436 393916 211488 393922
rect 211436 393858 211488 393864
rect 211448 14550 211476 393858
rect 211620 393848 211672 393854
rect 211620 393790 211672 393796
rect 211528 177336 211580 177342
rect 211528 177278 211580 177284
rect 211436 14544 211488 14550
rect 211436 14486 211488 14492
rect 211344 14476 211396 14482
rect 211344 14418 211396 14424
rect 210240 13184 210292 13190
rect 210240 13126 210292 13132
rect 210148 13116 210200 13122
rect 210148 13058 210200 13064
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 210056 9036 210108 9042
rect 210056 8978 210108 8984
rect 209964 8968 210016 8974
rect 209964 8910 210016 8916
rect 209792 6886 209912 6914
rect 209044 3868 209096 3874
rect 209044 3810 209096 3816
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 211540 6914 211568 177278
rect 211632 11830 211660 393790
rect 211816 14618 211844 397559
rect 211908 178702 211936 398550
rect 212000 394398 212028 400044
rect 211988 394392 212040 394398
rect 211988 394334 212040 394340
rect 212092 393922 212120 400044
rect 212184 397662 212212 400044
rect 212276 397730 212304 400044
rect 212264 397724 212316 397730
rect 212264 397666 212316 397672
rect 212172 397656 212224 397662
rect 212172 397598 212224 397604
rect 212172 397520 212224 397526
rect 212172 397462 212224 397468
rect 212080 393916 212132 393922
rect 212080 393858 212132 393864
rect 212184 393802 212212 397462
rect 212368 393854 212396 400044
rect 212460 398138 212488 400044
rect 212448 398132 212500 398138
rect 212448 398074 212500 398080
rect 212446 398032 212502 398041
rect 212446 397967 212502 397976
rect 212000 393774 212212 393802
rect 212356 393848 212408 393854
rect 212356 393790 212408 393796
rect 212000 354142 212028 393774
rect 212460 393666 212488 397967
rect 212552 397769 212580 400044
rect 212538 397760 212594 397769
rect 212538 397695 212594 397704
rect 212644 397497 212672 400044
rect 212630 397488 212686 397497
rect 212630 397423 212686 397432
rect 212736 395418 212764 400044
rect 212828 398449 212856 400044
rect 212814 398440 212870 398449
rect 212814 398375 212870 398384
rect 212816 397996 212868 398002
rect 212816 397938 212868 397944
rect 212828 397526 212856 397938
rect 212816 397520 212868 397526
rect 212816 397462 212868 397468
rect 212724 395412 212776 395418
rect 212724 395354 212776 395360
rect 212540 394392 212592 394398
rect 212540 394334 212592 394340
rect 212092 393638 212488 393666
rect 212092 354210 212120 393638
rect 212552 393530 212580 394334
rect 212920 394040 212948 400044
rect 213012 397633 213040 400044
rect 212998 397624 213054 397633
rect 212998 397559 213054 397568
rect 212736 394012 212948 394040
rect 212632 393984 212684 393990
rect 212632 393926 212684 393932
rect 212460 393502 212580 393530
rect 212460 389174 212488 393502
rect 212368 389146 212488 389174
rect 212080 354204 212132 354210
rect 212080 354146 212132 354152
rect 211988 354136 212040 354142
rect 211988 354078 212040 354084
rect 211896 178696 211948 178702
rect 211896 178638 211948 178644
rect 211804 14612 211856 14618
rect 211804 14554 211856 14560
rect 211620 11824 211672 11830
rect 211620 11766 211672 11772
rect 212368 11762 212396 389146
rect 212644 11966 212672 393926
rect 212632 11960 212684 11966
rect 212632 11902 212684 11908
rect 212736 11898 212764 394012
rect 213104 393938 213132 400044
rect 213196 393990 213224 400044
rect 212816 393916 212868 393922
rect 212816 393858 212868 393864
rect 212920 393910 213132 393938
rect 213184 393984 213236 393990
rect 213184 393926 213236 393932
rect 212828 14686 212856 393858
rect 212920 15910 212948 393910
rect 213288 393802 213316 400044
rect 213380 398177 213408 400044
rect 213366 398168 213422 398177
rect 213366 398103 213422 398112
rect 213368 397656 213420 397662
rect 213368 397598 213420 397604
rect 213012 393774 213316 393802
rect 213012 355366 213040 393774
rect 213092 393712 213144 393718
rect 213092 393654 213144 393660
rect 213104 355434 213132 393654
rect 213380 393394 213408 397598
rect 213472 396710 213500 400044
rect 213564 398614 213592 400044
rect 213552 398608 213604 398614
rect 213552 398550 213604 398556
rect 213460 396704 213512 396710
rect 213460 396646 213512 396652
rect 213656 393718 213684 400044
rect 213644 393712 213696 393718
rect 213644 393654 213696 393660
rect 213196 393366 213408 393394
rect 213092 355428 213144 355434
rect 213092 355370 213144 355376
rect 213000 355360 213052 355366
rect 213000 355302 213052 355308
rect 213196 354414 213224 393366
rect 213748 389174 213776 400044
rect 213840 393922 213868 400044
rect 213932 399129 213960 400044
rect 213918 399120 213974 399129
rect 213918 399055 213974 399064
rect 214024 398970 214052 400044
rect 213932 398942 214052 398970
rect 213932 397905 213960 398942
rect 214010 398032 214066 398041
rect 214010 397967 214066 397976
rect 213918 397896 213974 397905
rect 213918 397831 213974 397840
rect 213920 397724 213972 397730
rect 213920 397666 213972 397672
rect 213932 396914 213960 397666
rect 214024 397633 214052 397967
rect 214010 397624 214066 397633
rect 214010 397559 214066 397568
rect 214116 397497 214144 400044
rect 214208 397633 214236 400044
rect 214300 397769 214328 400044
rect 214286 397760 214342 397769
rect 214286 397695 214342 397704
rect 214194 397624 214250 397633
rect 214194 397559 214250 397568
rect 214102 397488 214158 397497
rect 214102 397423 214158 397432
rect 213920 396908 213972 396914
rect 213920 396850 213972 396856
rect 214392 394482 214420 400044
rect 214484 398993 214512 400044
rect 214470 398984 214526 398993
rect 214470 398919 214526 398928
rect 214470 398848 214526 398857
rect 214470 398783 214526 398792
rect 214484 395486 214512 398783
rect 214472 395480 214524 395486
rect 214472 395422 214524 395428
rect 214208 394454 214420 394482
rect 214012 393984 214064 393990
rect 214012 393926 214064 393932
rect 213828 393916 213880 393922
rect 213828 393858 213880 393864
rect 213288 389146 213776 389174
rect 213184 354408 213236 354414
rect 213184 354350 213236 354356
rect 212908 15904 212960 15910
rect 212908 15846 212960 15852
rect 212816 14680 212868 14686
rect 212816 14622 212868 14628
rect 213288 12034 213316 389146
rect 213276 12028 213328 12034
rect 213276 11970 213328 11976
rect 212724 11892 212776 11898
rect 212724 11834 212776 11840
rect 212356 11756 212408 11762
rect 212356 11698 212408 11704
rect 214024 9110 214052 393926
rect 214104 393780 214156 393786
rect 214104 393722 214156 393728
rect 214116 9178 214144 393722
rect 214208 12102 214236 394454
rect 214288 394392 214340 394398
rect 214576 394346 214604 400044
rect 214668 394398 214696 400044
rect 214288 394334 214340 394340
rect 214300 13258 214328 394334
rect 214484 394318 214604 394346
rect 214656 394392 214708 394398
rect 214656 394334 214708 394340
rect 214484 394040 214512 394318
rect 214484 394012 214696 394040
rect 214564 393916 214616 393922
rect 214564 393858 214616 393864
rect 214380 393848 214432 393854
rect 214380 393790 214432 393796
rect 214392 13326 214420 393790
rect 214472 390448 214524 390454
rect 214472 390390 214524 390396
rect 214484 354006 214512 390390
rect 214576 354074 214604 393858
rect 214668 389174 214696 394012
rect 214760 390454 214788 400044
rect 214852 393990 214880 400044
rect 214840 393984 214892 393990
rect 214840 393926 214892 393932
rect 214944 393854 214972 400044
rect 215036 397594 215064 400044
rect 215024 397588 215076 397594
rect 215024 397530 215076 397536
rect 214932 393848 214984 393854
rect 214932 393790 214984 393796
rect 215128 393786 215156 400044
rect 215220 393922 215248 400044
rect 215312 397497 215340 400044
rect 215298 397488 215354 397497
rect 215298 397423 215354 397432
rect 215404 396681 215432 400044
rect 215496 397633 215524 400044
rect 215588 397769 215616 400044
rect 215574 397760 215630 397769
rect 215574 397695 215630 397704
rect 215482 397624 215538 397633
rect 215482 397559 215538 397568
rect 215390 396672 215446 396681
rect 215390 396607 215446 396616
rect 215300 394528 215352 394534
rect 215300 394470 215352 394476
rect 215312 394194 215340 394470
rect 215300 394188 215352 394194
rect 215300 394130 215352 394136
rect 215680 394126 215708 400044
rect 215668 394120 215720 394126
rect 215668 394062 215720 394068
rect 215576 394052 215628 394058
rect 215576 393994 215628 394000
rect 215208 393916 215260 393922
rect 215208 393858 215260 393864
rect 215484 393916 215536 393922
rect 215484 393858 215536 393864
rect 215116 393780 215168 393786
rect 215116 393722 215168 393728
rect 214748 390448 214800 390454
rect 214748 390390 214800 390396
rect 214668 389146 214788 389174
rect 214564 354068 214616 354074
rect 214564 354010 214616 354016
rect 214472 354000 214524 354006
rect 214472 353942 214524 353948
rect 214380 13320 214432 13326
rect 214380 13262 214432 13268
rect 214288 13252 214340 13258
rect 214288 13194 214340 13200
rect 214196 12096 214248 12102
rect 214196 12038 214248 12044
rect 214104 9172 214156 9178
rect 214104 9114 214156 9120
rect 214012 9104 214064 9110
rect 214012 9046 214064 9052
rect 214760 7614 214788 389146
rect 215496 9314 215524 393858
rect 215588 13530 215616 393994
rect 215668 393984 215720 393990
rect 215668 393926 215720 393932
rect 215576 13524 215628 13530
rect 215576 13466 215628 13472
rect 215680 13462 215708 393926
rect 215668 13456 215720 13462
rect 215668 13398 215720 13404
rect 215772 13394 215800 400044
rect 215864 398177 215892 400044
rect 215850 398168 215906 398177
rect 215850 398103 215906 398112
rect 215956 393972 215984 400044
rect 216048 393990 216076 400044
rect 215864 393944 215984 393972
rect 216036 393984 216088 393990
rect 215864 391678 215892 393944
rect 216036 393926 216088 393932
rect 216140 391898 216168 400044
rect 216232 393922 216260 400044
rect 216324 394058 216352 400044
rect 216416 397730 216444 400044
rect 216404 397724 216456 397730
rect 216404 397666 216456 397672
rect 216404 397588 216456 397594
rect 216404 397530 216456 397536
rect 216312 394052 216364 394058
rect 216312 393994 216364 394000
rect 216220 393916 216272 393922
rect 216220 393858 216272 393864
rect 215956 391870 216168 391898
rect 216416 391882 216444 397530
rect 216404 391876 216456 391882
rect 215852 391672 215904 391678
rect 215852 391614 215904 391620
rect 215852 391536 215904 391542
rect 215852 391478 215904 391484
rect 215864 13598 215892 391478
rect 215956 14754 215984 391870
rect 216404 391818 216456 391824
rect 216036 391808 216088 391814
rect 216508 391762 216536 400044
rect 216036 391750 216088 391756
rect 216048 177546 216076 391750
rect 216140 391734 216536 391762
rect 216036 177540 216088 177546
rect 216036 177482 216088 177488
rect 215944 14748 215996 14754
rect 215944 14690 215996 14696
rect 215852 13592 215904 13598
rect 215852 13534 215904 13540
rect 215760 13388 215812 13394
rect 215760 13330 215812 13336
rect 216140 9382 216168 391734
rect 216220 391672 216272 391678
rect 216220 391614 216272 391620
rect 216128 9376 216180 9382
rect 216128 9318 216180 9324
rect 215484 9308 215536 9314
rect 215484 9250 215536 9256
rect 216232 9246 216260 391614
rect 216600 391542 216628 400044
rect 216692 397769 216720 400044
rect 216678 397760 216734 397769
rect 216678 397695 216734 397704
rect 216784 397497 216812 400044
rect 216876 397633 216904 400044
rect 216968 399265 216996 400044
rect 216954 399256 217010 399265
rect 216954 399191 217010 399200
rect 216956 399084 217008 399090
rect 216956 399026 217008 399032
rect 216862 397624 216918 397633
rect 216862 397559 216918 397568
rect 216770 397488 216826 397497
rect 216770 397423 216826 397432
rect 216968 395622 216996 399026
rect 217060 397905 217088 400044
rect 217046 397896 217102 397905
rect 217046 397831 217102 397840
rect 216956 395616 217008 395622
rect 216956 395558 217008 395564
rect 217048 394120 217100 394126
rect 217048 394062 217100 394068
rect 216956 394052 217008 394058
rect 216956 393994 217008 394000
rect 216864 393984 216916 393990
rect 216864 393926 216916 393932
rect 216772 393916 216824 393922
rect 216772 393858 216824 393864
rect 216588 391536 216640 391542
rect 216588 391478 216640 391484
rect 216784 10538 216812 393858
rect 216772 10532 216824 10538
rect 216772 10474 216824 10480
rect 216876 10470 216904 393926
rect 216968 14822 216996 393994
rect 217060 354346 217088 394062
rect 217048 354340 217100 354346
rect 217048 354282 217100 354288
rect 217152 354278 217180 400044
rect 217244 397662 217272 400044
rect 217232 397656 217284 397662
rect 217232 397598 217284 397604
rect 217336 393972 217364 400044
rect 217428 394126 217456 400044
rect 217416 394120 217468 394126
rect 217416 394062 217468 394068
rect 217336 393944 217456 393972
rect 217232 390312 217284 390318
rect 217232 390254 217284 390260
rect 217244 355502 217272 390254
rect 217232 355496 217284 355502
rect 217232 355438 217284 355444
rect 217140 354272 217192 354278
rect 217140 354214 217192 354220
rect 217048 177540 217100 177546
rect 217048 177482 217100 177488
rect 216956 14816 217008 14822
rect 216956 14758 217008 14764
rect 216864 10464 216916 10470
rect 216864 10406 216916 10412
rect 216220 9240 216272 9246
rect 216220 9182 216272 9188
rect 214748 7608 214800 7614
rect 214748 7550 214800 7556
rect 211540 6886 211752 6914
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 6886
rect 215668 3800 215720 3806
rect 215668 3742 215720 3748
rect 214472 3732 214524 3738
rect 214472 3674 214524 3680
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 213380 480 213408 3606
rect 214484 480 214512 3674
rect 215680 480 215708 3742
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 354 216946 480
rect 217060 354 217088 177482
rect 217428 10402 217456 393944
rect 217520 390318 217548 400044
rect 217612 393990 217640 400044
rect 217704 399090 217732 400044
rect 217692 399084 217744 399090
rect 217692 399026 217744 399032
rect 217692 398744 217744 398750
rect 217692 398686 217744 398692
rect 217600 393984 217652 393990
rect 217600 393926 217652 393932
rect 217508 390312 217560 390318
rect 217508 390254 217560 390260
rect 217704 389174 217732 398686
rect 217796 397934 217824 400044
rect 217784 397928 217836 397934
rect 217784 397870 217836 397876
rect 217784 397724 217836 397730
rect 217784 397666 217836 397672
rect 217796 392698 217824 397666
rect 217888 393922 217916 400044
rect 217980 394058 218008 400044
rect 218072 397497 218100 400044
rect 218058 397488 218114 397497
rect 218058 397423 218114 397432
rect 218164 396817 218192 400044
rect 218256 397633 218284 400044
rect 218348 397798 218376 400044
rect 218336 397792 218388 397798
rect 218336 397734 218388 397740
rect 218242 397624 218298 397633
rect 218242 397559 218298 397568
rect 218150 396808 218206 396817
rect 218150 396743 218206 396752
rect 218440 394074 218468 400044
rect 217968 394052 218020 394058
rect 217968 393994 218020 394000
rect 218256 394046 218468 394074
rect 217876 393916 217928 393922
rect 217876 393858 217928 393864
rect 217784 392692 217836 392698
rect 217784 392634 217836 392640
rect 217704 389146 218008 389174
rect 217416 10396 217468 10402
rect 217416 10338 217468 10344
rect 217980 4078 218008 389146
rect 218256 10606 218284 394046
rect 218532 393972 218560 400044
rect 218624 398138 218652 400044
rect 218612 398132 218664 398138
rect 218612 398074 218664 398080
rect 218440 393944 218560 393972
rect 218612 393984 218664 393990
rect 218336 393916 218388 393922
rect 218336 393858 218388 393864
rect 218348 10810 218376 393858
rect 218440 14890 218468 393944
rect 218612 393926 218664 393932
rect 218520 393848 218572 393854
rect 218520 393790 218572 393796
rect 218532 15978 218560 393790
rect 218624 354482 218652 393926
rect 218716 392562 218744 400044
rect 218808 394074 218836 400044
rect 218900 398478 218928 400044
rect 218888 398472 218940 398478
rect 218888 398414 218940 398420
rect 218888 398200 218940 398206
rect 218888 398142 218940 398148
rect 218900 395554 218928 398142
rect 218888 395548 218940 395554
rect 218888 395490 218940 395496
rect 218808 394046 218928 394074
rect 218900 392630 218928 394046
rect 218888 392624 218940 392630
rect 218888 392566 218940 392572
rect 218704 392556 218756 392562
rect 218704 392498 218756 392504
rect 218992 392442 219020 400044
rect 219084 393990 219112 400044
rect 219072 393984 219124 393990
rect 219072 393926 219124 393932
rect 219176 393854 219204 400044
rect 219268 393922 219296 400044
rect 219360 398206 219388 400044
rect 219452 398818 219480 400044
rect 219440 398812 219492 398818
rect 219440 398754 219492 398760
rect 219348 398200 219400 398206
rect 219348 398142 219400 398148
rect 219348 398064 219400 398070
rect 219348 398006 219400 398012
rect 219256 393916 219308 393922
rect 219256 393858 219308 393864
rect 219164 393848 219216 393854
rect 219164 393790 219216 393796
rect 218716 392414 219020 392442
rect 218612 354476 218664 354482
rect 218612 354418 218664 354424
rect 218612 46368 218664 46374
rect 218612 46310 218664 46316
rect 218520 15972 218572 15978
rect 218520 15914 218572 15920
rect 218428 14884 218480 14890
rect 218428 14826 218480 14832
rect 218336 10804 218388 10810
rect 218336 10746 218388 10752
rect 218244 10600 218296 10606
rect 218244 10542 218296 10548
rect 218624 6914 218652 46310
rect 218716 10742 218744 392414
rect 218796 392352 218848 392358
rect 218796 392294 218848 392300
rect 218704 10736 218756 10742
rect 218704 10678 218756 10684
rect 218808 10674 218836 392294
rect 218796 10668 218848 10674
rect 218796 10610 218848 10616
rect 218072 6886 218652 6914
rect 217968 4072 218020 4078
rect 217968 4014 218020 4020
rect 218072 480 218100 6886
rect 219256 4004 219308 4010
rect 219256 3946 219308 3952
rect 219268 480 219296 3946
rect 219360 3874 219388 398006
rect 219440 397724 219492 397730
rect 219440 397666 219492 397672
rect 219348 3868 219400 3874
rect 219348 3810 219400 3816
rect 219452 490 219480 397666
rect 219544 397497 219572 400044
rect 219530 397488 219586 397497
rect 219530 397423 219586 397432
rect 219636 395729 219664 400044
rect 219728 397497 219756 400044
rect 219820 397633 219848 400044
rect 219806 397624 219862 397633
rect 219806 397559 219862 397568
rect 219714 397488 219770 397497
rect 219714 397423 219770 397432
rect 219622 395720 219678 395729
rect 219622 395655 219678 395664
rect 219532 394120 219584 394126
rect 219532 394062 219584 394068
rect 219544 3602 219572 394062
rect 219624 394052 219676 394058
rect 219624 393994 219676 394000
rect 219532 3596 219584 3602
rect 219532 3538 219584 3544
rect 219636 3534 219664 393994
rect 219808 393984 219860 393990
rect 219912 393972 219940 400044
rect 220004 394074 220032 400044
rect 220096 397526 220124 400044
rect 220084 397520 220136 397526
rect 220084 397462 220136 397468
rect 220004 394046 220124 394074
rect 220188 394058 220216 400044
rect 219912 393944 220032 393972
rect 219808 393926 219860 393932
rect 219716 393916 219768 393922
rect 219716 393858 219768 393864
rect 219728 4894 219756 393858
rect 219820 6186 219848 393926
rect 219900 393848 219952 393854
rect 219900 393790 219952 393796
rect 219912 6254 219940 393790
rect 220004 14958 220032 393944
rect 220096 177410 220124 394046
rect 220176 394052 220228 394058
rect 220176 393994 220228 394000
rect 220280 393990 220308 400044
rect 220372 394126 220400 400044
rect 220464 394194 220492 400044
rect 220556 396846 220584 400044
rect 220544 396840 220596 396846
rect 220544 396782 220596 396788
rect 220452 394188 220504 394194
rect 220452 394130 220504 394136
rect 220360 394120 220412 394126
rect 220360 394062 220412 394068
rect 220268 393984 220320 393990
rect 220268 393926 220320 393932
rect 220648 393922 220676 400044
rect 220636 393916 220688 393922
rect 220636 393858 220688 393864
rect 220740 393854 220768 400044
rect 220832 399022 220860 400044
rect 220820 399016 220872 399022
rect 220820 398958 220872 398964
rect 220924 397633 220952 400044
rect 220910 397624 220966 397633
rect 220910 397559 220966 397568
rect 221016 397497 221044 400044
rect 221108 397633 221136 400044
rect 221094 397624 221150 397633
rect 221094 397559 221150 397568
rect 221200 397497 221228 400044
rect 221002 397488 221058 397497
rect 221002 397423 221058 397432
rect 221186 397488 221242 397497
rect 221186 397423 221242 397432
rect 221292 394330 221320 400044
rect 221280 394324 221332 394330
rect 221280 394266 221332 394272
rect 221004 394188 221056 394194
rect 221004 394130 221056 394136
rect 220912 394052 220964 394058
rect 220912 393994 220964 394000
rect 220728 393848 220780 393854
rect 220728 393790 220780 393796
rect 220084 177404 220136 177410
rect 220084 177346 220136 177352
rect 219992 14952 220044 14958
rect 219992 14894 220044 14900
rect 219900 6248 219952 6254
rect 219900 6190 219952 6196
rect 219808 6180 219860 6186
rect 219808 6122 219860 6128
rect 220924 5030 220952 393994
rect 220912 5024 220964 5030
rect 220912 4966 220964 4972
rect 221016 4962 221044 394130
rect 221188 394120 221240 394126
rect 221188 394062 221240 394068
rect 221096 393984 221148 393990
rect 221096 393926 221148 393932
rect 221108 7886 221136 393926
rect 221200 393904 221228 394062
rect 221200 393876 221320 393904
rect 221188 393780 221240 393786
rect 221188 393722 221240 393728
rect 221096 7880 221148 7886
rect 221096 7822 221148 7828
rect 221200 7818 221228 393722
rect 221188 7812 221240 7818
rect 221188 7754 221240 7760
rect 221292 7750 221320 393876
rect 221280 7744 221332 7750
rect 221280 7686 221332 7692
rect 221384 7682 221412 400044
rect 221476 394194 221504 400044
rect 221464 394188 221516 394194
rect 221464 394130 221516 394136
rect 221568 394126 221596 400044
rect 221660 397050 221688 400044
rect 221648 397044 221700 397050
rect 221648 396986 221700 396992
rect 221648 394324 221700 394330
rect 221648 394266 221700 394272
rect 221556 394120 221608 394126
rect 221556 394062 221608 394068
rect 221660 393972 221688 394266
rect 221752 394058 221780 400044
rect 221740 394052 221792 394058
rect 221740 393994 221792 394000
rect 221568 393944 221688 393972
rect 221464 393236 221516 393242
rect 221464 393178 221516 393184
rect 221476 46238 221504 393178
rect 221568 177478 221596 393944
rect 221844 393786 221872 400044
rect 221832 393780 221884 393786
rect 221832 393722 221884 393728
rect 221936 393242 221964 400044
rect 221924 393236 221976 393242
rect 221924 393178 221976 393184
rect 222028 389174 222056 400044
rect 222120 393990 222148 400044
rect 222212 397769 222240 400044
rect 222198 397760 222254 397769
rect 222198 397695 222254 397704
rect 222200 397656 222252 397662
rect 222200 397598 222252 397604
rect 222108 393984 222160 393990
rect 222108 393926 222160 393932
rect 221660 389146 222056 389174
rect 221556 177472 221608 177478
rect 221556 177414 221608 177420
rect 221464 46232 221516 46238
rect 221464 46174 221516 46180
rect 221372 7676 221424 7682
rect 221372 7618 221424 7624
rect 221660 5098 221688 389146
rect 222212 16574 222240 397598
rect 222304 397497 222332 400044
rect 222396 397594 222424 400044
rect 222384 397588 222436 397594
rect 222384 397530 222436 397536
rect 222290 397488 222346 397497
rect 222290 397423 222346 397432
rect 222488 397118 222516 400044
rect 222476 397112 222528 397118
rect 222476 397054 222528 397060
rect 222384 394052 222436 394058
rect 222384 393994 222436 394000
rect 222212 16546 222332 16574
rect 221648 5092 221700 5098
rect 221648 5034 221700 5040
rect 221004 4956 221056 4962
rect 221004 4898 221056 4904
rect 219716 4888 219768 4894
rect 219716 4830 219768 4836
rect 219624 3528 219676 3534
rect 219624 3470 219676 3476
rect 222304 3482 222332 16546
rect 222396 5302 222424 393994
rect 222476 393984 222528 393990
rect 222476 393926 222528 393932
rect 222384 5296 222436 5302
rect 222384 5238 222436 5244
rect 222488 5234 222516 393926
rect 222580 390046 222608 400044
rect 222568 390040 222620 390046
rect 222568 389982 222620 389988
rect 222568 389904 222620 389910
rect 222568 389846 222620 389852
rect 222580 6322 222608 389846
rect 222672 7954 222700 400044
rect 222764 393922 222792 400044
rect 222856 397798 222884 400044
rect 222844 397792 222896 397798
rect 222844 397734 222896 397740
rect 222948 393990 222976 400044
rect 222936 393984 222988 393990
rect 222936 393926 222988 393932
rect 222752 393916 222804 393922
rect 222752 393858 222804 393864
rect 223040 393768 223068 400044
rect 223132 398002 223160 400044
rect 223120 397996 223172 398002
rect 223120 397938 223172 397944
rect 223120 395548 223172 395554
rect 223120 395490 223172 395496
rect 222764 393740 223068 393768
rect 222764 46306 222792 393740
rect 223132 392442 223160 395490
rect 223224 394058 223252 400044
rect 223212 394052 223264 394058
rect 223212 393994 223264 394000
rect 223212 393916 223264 393922
rect 223212 393858 223264 393864
rect 222856 392414 223160 392442
rect 222752 46300 222804 46306
rect 222752 46242 222804 46248
rect 222660 7948 222712 7954
rect 222660 7890 222712 7896
rect 222568 6316 222620 6322
rect 222568 6258 222620 6264
rect 222476 5228 222528 5234
rect 222476 5170 222528 5176
rect 222856 4010 222884 392414
rect 222936 392216 222988 392222
rect 223224 392170 223252 393858
rect 223316 392222 223344 400044
rect 223408 398682 223436 400044
rect 223396 398676 223448 398682
rect 223396 398618 223448 398624
rect 222936 392158 222988 392164
rect 222948 177614 222976 392158
rect 223040 392142 223252 392170
rect 223304 392216 223356 392222
rect 223304 392158 223356 392164
rect 223040 352646 223068 392142
rect 223212 390040 223264 390046
rect 223212 389982 223264 389988
rect 223028 352640 223080 352646
rect 223028 352582 223080 352588
rect 222936 177608 222988 177614
rect 222936 177550 222988 177556
rect 223224 5166 223252 389982
rect 223500 389910 223528 400044
rect 223592 397905 223620 400044
rect 223684 398274 223712 400044
rect 223672 398268 223724 398274
rect 223672 398210 223724 398216
rect 223578 397896 223634 397905
rect 223578 397831 223634 397840
rect 223776 397497 223804 400044
rect 223868 397769 223896 400044
rect 223854 397760 223910 397769
rect 223854 397695 223910 397704
rect 223960 397633 223988 400044
rect 223946 397624 224002 397633
rect 223946 397559 224002 397568
rect 223762 397488 223818 397497
rect 223762 397423 223818 397432
rect 223672 394052 223724 394058
rect 223672 393994 223724 394000
rect 223488 389904 223540 389910
rect 223488 389846 223540 389852
rect 223212 5160 223264 5166
rect 223212 5102 223264 5108
rect 222844 4004 222896 4010
rect 222844 3946 222896 3952
rect 222304 3454 222792 3482
rect 223684 3466 223712 393994
rect 223856 393984 223908 393990
rect 224052 393972 224080 400044
rect 223856 393926 223908 393932
rect 223960 393944 224080 393972
rect 223764 389836 223816 389842
rect 223764 389778 223816 389784
rect 223776 6526 223804 389778
rect 223868 6594 223896 393926
rect 223856 6588 223908 6594
rect 223856 6530 223908 6536
rect 223764 6520 223816 6526
rect 223764 6462 223816 6468
rect 223960 6390 223988 393944
rect 224040 393848 224092 393854
rect 224040 393790 224092 393796
rect 224052 6458 224080 393790
rect 224144 178770 224172 400044
rect 224236 394534 224264 400044
rect 224224 394528 224276 394534
rect 224224 394470 224276 394476
rect 224328 393854 224356 400044
rect 224316 393848 224368 393854
rect 224316 393790 224368 393796
rect 224420 393666 224448 400044
rect 224512 394058 224540 400044
rect 224500 394052 224552 394058
rect 224500 393994 224552 394000
rect 224236 393638 224448 393666
rect 224236 352714 224264 393638
rect 224604 389842 224632 400044
rect 224696 397254 224724 400044
rect 224684 397248 224736 397254
rect 224684 397190 224736 397196
rect 224592 389836 224644 389842
rect 224592 389778 224644 389784
rect 224788 389174 224816 400044
rect 224880 393990 224908 400044
rect 224972 397769 225000 400044
rect 225064 398342 225092 400044
rect 225052 398336 225104 398342
rect 225052 398278 225104 398284
rect 224958 397760 225014 397769
rect 224958 397695 225014 397704
rect 225156 397497 225184 400044
rect 225248 397633 225276 400044
rect 225234 397624 225290 397633
rect 225234 397559 225290 397568
rect 225142 397488 225198 397497
rect 225142 397423 225198 397432
rect 225340 397066 225368 400044
rect 225432 397905 225460 400044
rect 225418 397896 225474 397905
rect 225418 397831 225474 397840
rect 225524 397186 225552 400044
rect 225512 397180 225564 397186
rect 225512 397122 225564 397128
rect 225616 397118 225644 400044
rect 225064 397038 225368 397066
rect 225604 397112 225656 397118
rect 225604 397054 225656 397060
rect 225064 394330 225092 397038
rect 225328 396908 225380 396914
rect 225708 396896 225736 400044
rect 225328 396850 225380 396856
rect 225432 396868 225736 396896
rect 225144 396704 225196 396710
rect 225144 396646 225196 396652
rect 225052 394324 225104 394330
rect 225052 394266 225104 394272
rect 224868 393984 224920 393990
rect 224868 393926 224920 393932
rect 224328 389146 224816 389174
rect 224224 352708 224276 352714
rect 224224 352650 224276 352656
rect 224132 178764 224184 178770
rect 224132 178706 224184 178712
rect 224040 6452 224092 6458
rect 224040 6394 224092 6400
rect 223948 6384 224000 6390
rect 223948 6326 224000 6332
rect 223948 4072 224000 4078
rect 223948 4014 224000 4020
rect 221556 3392 221608 3398
rect 221556 3334 221608 3340
rect 216834 326 217088 354
rect 216834 -960 216946 326
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 219452 462 220032 490
rect 221568 480 221596 3334
rect 222764 480 222792 3454
rect 223672 3460 223724 3466
rect 223672 3402 223724 3408
rect 223960 480 223988 4014
rect 224328 3942 224356 389146
rect 225156 4826 225184 396646
rect 225236 394596 225288 394602
rect 225236 394538 225288 394544
rect 225144 4820 225196 4826
rect 225144 4762 225196 4768
rect 224316 3936 224368 3942
rect 224316 3878 224368 3884
rect 225248 1578 225276 394538
rect 225340 6662 225368 396850
rect 225432 8022 225460 396868
rect 225800 396794 225828 400044
rect 225892 396914 225920 400044
rect 225880 396908 225932 396914
rect 225880 396850 225932 396856
rect 225524 396766 225828 396794
rect 225524 352782 225552 396766
rect 225984 396642 226012 400044
rect 226076 397322 226104 400044
rect 226064 397316 226116 397322
rect 226064 397258 226116 397264
rect 226064 397112 226116 397118
rect 226064 397054 226116 397060
rect 225788 396636 225840 396642
rect 225788 396578 225840 396584
rect 225972 396636 226024 396642
rect 225972 396578 226024 396584
rect 225604 396568 225656 396574
rect 225604 396510 225656 396516
rect 225512 352776 225564 352782
rect 225512 352718 225564 352724
rect 225420 8016 225472 8022
rect 225420 7958 225472 7964
rect 225328 6656 225380 6662
rect 225328 6598 225380 6604
rect 225616 3806 225644 396510
rect 225696 351960 225748 351966
rect 225696 351902 225748 351908
rect 225604 3800 225656 3806
rect 225604 3742 225656 3748
rect 225708 3398 225736 351902
rect 225800 5438 225828 396578
rect 226076 393314 226104 397054
rect 226168 394466 226196 400044
rect 226260 396710 226288 400044
rect 226352 398886 226380 400044
rect 226340 398880 226392 398886
rect 226340 398822 226392 398828
rect 226444 398410 226472 400044
rect 226536 398546 226564 400044
rect 226524 398540 226576 398546
rect 226524 398482 226576 398488
rect 226432 398404 226484 398410
rect 226432 398346 226484 398352
rect 226628 397610 226656 400044
rect 226720 398954 226748 400044
rect 226708 398948 226760 398954
rect 226708 398890 226760 398896
rect 226340 397588 226392 397594
rect 226340 397530 226392 397536
rect 226444 397582 226656 397610
rect 226248 396704 226300 396710
rect 226248 396646 226300 396652
rect 226156 394460 226208 394466
rect 226156 394402 226208 394408
rect 225892 393286 226104 393314
rect 225788 5432 225840 5438
rect 225788 5374 225840 5380
rect 225892 5370 225920 393286
rect 225880 5364 225932 5370
rect 225880 5306 225932 5312
rect 225696 3392 225748 3398
rect 225696 3334 225748 3340
rect 225156 1550 225276 1578
rect 225156 480 225184 1550
rect 226352 480 226380 397530
rect 226444 396409 226472 397582
rect 226616 396772 226668 396778
rect 226616 396714 226668 396720
rect 226524 396636 226576 396642
rect 226524 396578 226576 396584
rect 226430 396400 226486 396409
rect 226430 396335 226486 396344
rect 226536 3738 226564 396578
rect 226628 46374 226656 396714
rect 226708 396704 226760 396710
rect 226708 396646 226760 396652
rect 226720 177546 226748 396646
rect 226708 177540 226760 177546
rect 226708 177482 226760 177488
rect 226812 177342 226840 400044
rect 226904 396386 226932 400044
rect 226996 396642 227024 400044
rect 226984 396636 227036 396642
rect 226984 396578 227036 396584
rect 227088 396574 227116 400044
rect 227180 396710 227208 400044
rect 227272 396778 227300 400044
rect 227260 396772 227312 396778
rect 227260 396714 227312 396720
rect 227168 396704 227220 396710
rect 227168 396646 227220 396652
rect 227076 396568 227128 396574
rect 227076 396510 227128 396516
rect 226904 396358 227300 396386
rect 226892 396296 226944 396302
rect 226892 396238 226944 396244
rect 226904 351966 226932 396238
rect 227272 393314 227300 396358
rect 227364 395554 227392 400044
rect 227456 397730 227484 400044
rect 227444 397724 227496 397730
rect 227444 397666 227496 397672
rect 227548 396302 227576 400044
rect 227640 397662 227668 400044
rect 227732 398750 227760 400044
rect 227720 398744 227772 398750
rect 227720 398686 227772 398692
rect 227628 397656 227680 397662
rect 227628 397598 227680 397604
rect 227628 397520 227680 397526
rect 227628 397462 227680 397468
rect 227536 396296 227588 396302
rect 227536 396238 227588 396244
rect 227352 395548 227404 395554
rect 227352 395490 227404 395496
rect 227272 393286 227484 393314
rect 226892 351960 226944 351966
rect 226892 351902 226944 351908
rect 226800 177336 226852 177342
rect 226800 177278 226852 177284
rect 226892 176724 226944 176730
rect 226892 176666 226944 176672
rect 226616 46368 226668 46374
rect 226616 46310 226668 46316
rect 226904 16574 226932 176666
rect 226904 16546 227392 16574
rect 226524 3732 226576 3738
rect 226524 3674 226576 3680
rect 227364 3482 227392 16546
rect 227456 3670 227484 393286
rect 227444 3664 227496 3670
rect 227444 3606 227496 3612
rect 227364 3454 227576 3482
rect 227548 480 227576 3454
rect 227640 2922 227668 397462
rect 227824 397066 227852 400044
rect 227916 397594 227944 400044
rect 227904 397588 227956 397594
rect 227904 397530 227956 397536
rect 227732 397038 227852 397066
rect 227732 394602 227760 397038
rect 227812 396976 227864 396982
rect 227812 396918 227864 396924
rect 227824 396250 227852 396918
rect 228008 396506 228036 400044
rect 228100 396846 228128 400044
rect 228088 396840 228140 396846
rect 228088 396782 228140 396788
rect 227996 396500 228048 396506
rect 227996 396442 228048 396448
rect 228192 396386 228220 400044
rect 228284 397526 228312 400044
rect 228272 397520 228324 397526
rect 228272 397462 228324 397468
rect 228376 396794 228404 400044
rect 228100 396358 228220 396386
rect 228284 396766 228404 396794
rect 227824 396222 228036 396250
rect 227720 394596 227772 394602
rect 227720 394538 227772 394544
rect 227904 393372 227956 393378
rect 227904 393314 227956 393320
rect 227916 4010 227944 393314
rect 227904 4004 227956 4010
rect 227904 3946 227956 3952
rect 228008 3942 228036 396222
rect 228100 4146 228128 396358
rect 228180 396296 228232 396302
rect 228180 396238 228232 396244
rect 228192 176730 228220 396238
rect 228284 394738 228312 396766
rect 228364 395412 228416 395418
rect 228364 395354 228416 395360
rect 228272 394732 228324 394738
rect 228272 394674 228324 394680
rect 228272 394596 228324 394602
rect 228272 394538 228324 394544
rect 228284 177342 228312 394538
rect 228376 354142 228404 395354
rect 228468 393378 228496 400044
rect 228560 395418 228588 400044
rect 228652 396982 228680 400044
rect 228640 396976 228692 396982
rect 228640 396918 228692 396924
rect 228640 396840 228692 396846
rect 228640 396782 228692 396788
rect 228548 395412 228600 395418
rect 228548 395354 228600 395360
rect 228456 393372 228508 393378
rect 228456 393314 228508 393320
rect 228652 393314 228680 396782
rect 228560 393286 228680 393314
rect 228744 393314 228772 400044
rect 228836 394602 228864 400044
rect 228928 397497 228956 400044
rect 229020 397905 229048 400044
rect 229006 397896 229062 397905
rect 229006 397831 229062 397840
rect 228914 397488 228970 397497
rect 228914 397423 228970 397432
rect 229112 396574 229140 400044
rect 229204 397050 229232 400044
rect 229192 397044 229244 397050
rect 229192 396986 229244 396992
rect 229296 396982 229324 400044
rect 229284 396976 229336 396982
rect 229284 396918 229336 396924
rect 229388 396914 229416 400044
rect 229376 396908 229428 396914
rect 229376 396850 229428 396856
rect 229480 396794 229508 400044
rect 229204 396766 229508 396794
rect 229100 396568 229152 396574
rect 229100 396510 229152 396516
rect 228824 394596 228876 394602
rect 228824 394538 228876 394544
rect 228744 393286 229048 393314
rect 228364 354136 228416 354142
rect 228364 354078 228416 354084
rect 228272 177336 228324 177342
rect 228272 177278 228324 177284
rect 228180 176724 228232 176730
rect 228180 176666 228232 176672
rect 228088 4140 228140 4146
rect 228088 4082 228140 4088
rect 227996 3936 228048 3942
rect 227996 3878 228048 3884
rect 227628 2916 227680 2922
rect 227628 2858 227680 2864
rect 220004 354 220032 462
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228560 354 228588 393286
rect 229020 3670 229048 393286
rect 229008 3664 229060 3670
rect 229008 3606 229060 3612
rect 229204 3466 229232 396766
rect 229284 396704 229336 396710
rect 229572 396658 229600 400044
rect 229284 396646 229336 396652
rect 229192 3460 229244 3466
rect 229192 3402 229244 3408
rect 229296 3330 229324 396646
rect 229388 396630 229600 396658
rect 229664 396658 229692 400044
rect 229756 396778 229784 400044
rect 229744 396772 229796 396778
rect 229744 396714 229796 396720
rect 229664 396630 229784 396658
rect 229388 3602 229416 396630
rect 229468 396568 229520 396574
rect 229468 396510 229520 396516
rect 229652 396568 229704 396574
rect 229652 396510 229704 396516
rect 229480 4962 229508 396510
rect 229560 394256 229612 394262
rect 229560 394198 229612 394204
rect 229468 4956 229520 4962
rect 229468 4898 229520 4904
rect 229572 4826 229600 394198
rect 229664 4894 229692 396510
rect 229756 354074 229784 396630
rect 229848 396574 229876 400044
rect 229836 396568 229888 396574
rect 229836 396510 229888 396516
rect 229940 394262 229968 400044
rect 230032 397497 230060 400044
rect 230124 397633 230152 400044
rect 230216 398041 230244 400044
rect 230308 398206 230336 400044
rect 230296 398200 230348 398206
rect 230296 398142 230348 398148
rect 230202 398032 230258 398041
rect 230202 397967 230258 397976
rect 230400 397769 230428 400044
rect 230386 397760 230442 397769
rect 230386 397695 230442 397704
rect 230110 397624 230166 397633
rect 230110 397559 230166 397568
rect 230018 397488 230074 397497
rect 230018 397423 230074 397432
rect 230492 397118 230520 400044
rect 230480 397112 230532 397118
rect 230480 397054 230532 397060
rect 230204 397044 230256 397050
rect 230204 396986 230256 396992
rect 230112 396976 230164 396982
rect 230112 396918 230164 396924
rect 230020 396908 230072 396914
rect 230020 396850 230072 396856
rect 229928 394256 229980 394262
rect 229928 394198 229980 394204
rect 230032 393314 230060 396850
rect 229848 393286 230060 393314
rect 229744 354068 229796 354074
rect 229744 354010 229796 354016
rect 229848 354006 229876 393286
rect 229836 354000 229888 354006
rect 229836 353942 229888 353948
rect 229652 4888 229704 4894
rect 229652 4830 229704 4836
rect 229560 4820 229612 4826
rect 229560 4762 229612 4768
rect 229836 4140 229888 4146
rect 229836 4082 229888 4088
rect 229376 3596 229428 3602
rect 229376 3538 229428 3544
rect 229284 3324 229336 3330
rect 229284 3266 229336 3272
rect 229848 480 229876 4082
rect 230124 3398 230152 396918
rect 230216 394262 230244 396986
rect 230584 396846 230612 400044
rect 230572 396840 230624 396846
rect 230572 396782 230624 396788
rect 230572 396704 230624 396710
rect 230572 396646 230624 396652
rect 230676 396658 230704 400044
rect 230768 396778 230796 400044
rect 230860 398818 230888 400044
rect 230848 398812 230900 398818
rect 230848 398754 230900 398760
rect 230756 396772 230808 396778
rect 230756 396714 230808 396720
rect 230204 394256 230256 394262
rect 230204 394198 230256 394204
rect 230584 4146 230612 396646
rect 230676 396630 230888 396658
rect 230756 396568 230808 396574
rect 230756 396510 230808 396516
rect 230664 396500 230716 396506
rect 230664 396442 230716 396448
rect 230676 6798 230704 396442
rect 230768 6866 230796 396510
rect 230756 6860 230808 6866
rect 230756 6802 230808 6808
rect 230664 6792 230716 6798
rect 230664 6734 230716 6740
rect 230860 6050 230888 396630
rect 230952 6118 230980 400044
rect 231044 396914 231072 400044
rect 231032 396908 231084 396914
rect 231032 396850 231084 396856
rect 231032 396772 231084 396778
rect 231032 396714 231084 396720
rect 231044 354346 231072 396714
rect 231136 396574 231164 400044
rect 231124 396568 231176 396574
rect 231124 396510 231176 396516
rect 231228 396506 231256 400044
rect 231216 396500 231268 396506
rect 231216 396442 231268 396448
rect 231320 395758 231348 400044
rect 231412 396710 231440 400044
rect 231504 397526 231532 400044
rect 231596 397769 231624 400044
rect 231582 397760 231638 397769
rect 231582 397695 231638 397704
rect 231492 397520 231544 397526
rect 231688 397497 231716 400044
rect 231780 397633 231808 400044
rect 231766 397624 231822 397633
rect 231766 397559 231822 397568
rect 231492 397462 231544 397468
rect 231674 397488 231730 397497
rect 231674 397423 231730 397432
rect 231872 396982 231900 400044
rect 231964 397798 231992 400044
rect 231952 397792 232004 397798
rect 231952 397734 232004 397740
rect 231860 396976 231912 396982
rect 231860 396918 231912 396924
rect 231492 396908 231544 396914
rect 231492 396850 231544 396856
rect 231400 396704 231452 396710
rect 231400 396646 231452 396652
rect 231504 395826 231532 396850
rect 231768 396840 231820 396846
rect 231768 396782 231820 396788
rect 231860 396840 231912 396846
rect 231860 396782 231912 396788
rect 231492 395820 231544 395826
rect 231492 395762 231544 395768
rect 231308 395752 231360 395758
rect 231308 395694 231360 395700
rect 231124 394732 231176 394738
rect 231124 394674 231176 394680
rect 231032 354340 231084 354346
rect 231032 354282 231084 354288
rect 230940 6112 230992 6118
rect 230940 6054 230992 6060
rect 230848 6044 230900 6050
rect 230848 5986 230900 5992
rect 230572 4140 230624 4146
rect 230572 4082 230624 4088
rect 231136 3534 231164 394674
rect 231780 4078 231808 396782
rect 231872 17542 231900 396782
rect 232056 396658 232084 400044
rect 231964 396630 232084 396658
rect 232148 396658 232176 400044
rect 232240 396778 232268 400044
rect 232332 396846 232360 400044
rect 232320 396840 232372 396846
rect 232320 396782 232372 396788
rect 232228 396772 232280 396778
rect 232228 396714 232280 396720
rect 232424 396658 232452 400044
rect 232148 396630 232268 396658
rect 231964 17610 231992 396630
rect 232044 396568 232096 396574
rect 232044 396510 232096 396516
rect 232056 18970 232084 396510
rect 232136 396500 232188 396506
rect 232136 396442 232188 396448
rect 232148 25838 232176 396442
rect 232240 25974 232268 396630
rect 232332 396630 232452 396658
rect 232228 25968 232280 25974
rect 232228 25910 232280 25916
rect 232332 25906 232360 396630
rect 232412 394732 232464 394738
rect 232412 394674 232464 394680
rect 232424 87854 232452 394674
rect 232516 355502 232544 400044
rect 232608 396930 232636 400044
rect 232700 397050 232728 400044
rect 232688 397044 232740 397050
rect 232688 396986 232740 396992
rect 232608 396902 232728 396930
rect 232596 396772 232648 396778
rect 232596 396714 232648 396720
rect 232608 392766 232636 396714
rect 232700 396574 232728 396902
rect 232688 396568 232740 396574
rect 232688 396510 232740 396516
rect 232792 394738 232820 400044
rect 232884 397633 232912 400044
rect 232976 398041 233004 400044
rect 232962 398032 233018 398041
rect 232962 397967 233018 397976
rect 232870 397624 232926 397633
rect 232870 397559 232926 397568
rect 233068 397497 233096 400044
rect 233160 397769 233188 400044
rect 233252 398070 233280 400044
rect 233240 398064 233292 398070
rect 233240 398006 233292 398012
rect 233146 397760 233202 397769
rect 233146 397695 233202 397704
rect 233054 397488 233110 397497
rect 233054 397423 233110 397432
rect 232872 397044 232924 397050
rect 232872 396986 232924 396992
rect 232884 396506 232912 396986
rect 232964 396976 233016 396982
rect 232964 396918 233016 396924
rect 232872 396500 232924 396506
rect 232872 396442 232924 396448
rect 232976 395690 233004 396918
rect 232964 395684 233016 395690
rect 232964 395626 233016 395632
rect 232780 394732 232832 394738
rect 232780 394674 232832 394680
rect 232596 392760 232648 392766
rect 232596 392702 232648 392708
rect 232504 355496 232556 355502
rect 232504 355438 232556 355444
rect 232504 354136 232556 354142
rect 232504 354078 232556 354084
rect 232412 87848 232464 87854
rect 232412 87790 232464 87796
rect 232320 25900 232372 25906
rect 232320 25842 232372 25848
rect 232136 25832 232188 25838
rect 232136 25774 232188 25780
rect 232044 18964 232096 18970
rect 232044 18906 232096 18912
rect 231952 17604 232004 17610
rect 231952 17546 232004 17552
rect 231860 17536 231912 17542
rect 231860 17478 231912 17484
rect 231768 4072 231820 4078
rect 231768 4014 231820 4020
rect 231124 3528 231176 3534
rect 231124 3470 231176 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 230112 3392 230164 3398
rect 230112 3334 230164 3340
rect 231032 2916 231084 2922
rect 231032 2858 231084 2864
rect 231044 480 231072 2858
rect 232240 480 232268 3470
rect 232516 3126 232544 354078
rect 233344 3806 233372 400044
rect 233436 396658 233464 400044
rect 233528 396778 233556 400044
rect 233620 396846 233648 400044
rect 233608 396840 233660 396846
rect 233608 396782 233660 396788
rect 233516 396772 233568 396778
rect 233516 396714 233568 396720
rect 233436 396630 233648 396658
rect 233516 396568 233568 396574
rect 233516 396510 233568 396516
rect 233424 396500 233476 396506
rect 233424 396442 233476 396448
rect 233436 7818 233464 396442
rect 233528 18766 233556 396510
rect 233620 18902 233648 396630
rect 233608 18896 233660 18902
rect 233608 18838 233660 18844
rect 233712 18834 233740 400044
rect 233804 25770 233832 400044
rect 233896 398585 233924 400044
rect 233882 398576 233938 398585
rect 233882 398511 233938 398520
rect 233884 396772 233936 396778
rect 233884 396714 233936 396720
rect 233896 396386 233924 396714
rect 233988 396574 234016 400044
rect 234080 397662 234108 400044
rect 234068 397656 234120 397662
rect 234068 397598 234120 397604
rect 234068 397520 234120 397526
rect 234068 397462 234120 397468
rect 233976 396568 234028 396574
rect 233976 396510 234028 396516
rect 233896 396358 234016 396386
rect 233884 396296 233936 396302
rect 233884 396238 233936 396244
rect 233792 25764 233844 25770
rect 233792 25706 233844 25712
rect 233700 18828 233752 18834
rect 233700 18770 233752 18776
rect 233516 18760 233568 18766
rect 233516 18702 233568 18708
rect 233896 17678 233924 396238
rect 233988 389978 234016 396358
rect 234080 396302 234108 397462
rect 234172 396506 234200 400044
rect 234264 397497 234292 400044
rect 234356 397633 234384 400044
rect 234448 397769 234476 400044
rect 234434 397760 234490 397769
rect 234434 397695 234490 397704
rect 234436 397656 234488 397662
rect 234342 397624 234398 397633
rect 234436 397598 234488 397604
rect 234342 397559 234398 397568
rect 234250 397488 234306 397497
rect 234250 397423 234306 397432
rect 234252 396840 234304 396846
rect 234252 396782 234304 396788
rect 234160 396500 234212 396506
rect 234160 396442 234212 396448
rect 234068 396296 234120 396302
rect 234068 396238 234120 396244
rect 233976 389972 234028 389978
rect 233976 389914 234028 389920
rect 233884 17672 233936 17678
rect 233884 17614 233936 17620
rect 233424 7812 233476 7818
rect 233424 7754 233476 7760
rect 233424 4004 233476 4010
rect 233424 3946 233476 3952
rect 233332 3800 233384 3806
rect 233332 3742 233384 3748
rect 232504 3120 232556 3126
rect 232504 3062 232556 3068
rect 233436 480 233464 3946
rect 234264 3738 234292 396782
rect 234448 394534 234476 397598
rect 234540 397361 234568 400044
rect 234526 397352 234582 397361
rect 234526 397287 234582 397296
rect 234632 396930 234660 400044
rect 234724 397905 234752 400044
rect 234710 397896 234766 397905
rect 234710 397831 234766 397840
rect 234540 396902 234660 396930
rect 234540 396438 234568 396902
rect 234528 396432 234580 396438
rect 234528 396374 234580 396380
rect 234436 394528 234488 394534
rect 234436 394470 234488 394476
rect 234712 394392 234764 394398
rect 234712 394334 234764 394340
rect 234620 394120 234672 394126
rect 234620 394062 234672 394068
rect 234632 6730 234660 394062
rect 234724 7750 234752 394334
rect 234816 394040 234844 400044
rect 234908 394262 234936 400044
rect 234896 394256 234948 394262
rect 234896 394198 234948 394204
rect 235000 394126 235028 400044
rect 234988 394120 235040 394126
rect 234988 394062 235040 394068
rect 234816 394012 234936 394040
rect 234804 393848 234856 393854
rect 234804 393790 234856 393796
rect 234712 7744 234764 7750
rect 234712 7686 234764 7692
rect 234816 7682 234844 393790
rect 234908 18698 234936 394012
rect 234988 393984 235040 393990
rect 234988 393926 235040 393932
rect 235000 20262 235028 393926
rect 235092 20330 235120 400044
rect 235184 25702 235212 400044
rect 235276 394398 235304 400044
rect 235264 394392 235316 394398
rect 235264 394334 235316 394340
rect 235264 394256 235316 394262
rect 235264 394198 235316 394204
rect 235276 393836 235304 394198
rect 235368 393990 235396 400044
rect 235460 396658 235488 400044
rect 235552 396794 235580 400044
rect 235644 397225 235672 400044
rect 235736 397633 235764 400044
rect 235722 397624 235778 397633
rect 235722 397559 235778 397568
rect 235828 397497 235856 400044
rect 235920 397769 235948 400044
rect 235906 397760 235962 397769
rect 235906 397695 235962 397704
rect 235814 397488 235870 397497
rect 235814 397423 235870 397432
rect 235630 397216 235686 397225
rect 235630 397151 235686 397160
rect 235552 396766 235764 396794
rect 235460 396630 235580 396658
rect 235448 396432 235500 396438
rect 235448 396374 235500 396380
rect 235356 393984 235408 393990
rect 235356 393926 235408 393932
rect 235276 393808 235396 393836
rect 235264 393712 235316 393718
rect 235264 393654 235316 393660
rect 235276 87786 235304 393654
rect 235368 352714 235396 393808
rect 235460 393718 235488 396374
rect 235552 394466 235580 396630
rect 235540 394460 235592 394466
rect 235540 394402 235592 394408
rect 235736 393854 235764 396766
rect 236012 394670 236040 400044
rect 236104 397526 236132 400044
rect 236092 397520 236144 397526
rect 236092 397462 236144 397468
rect 236000 394664 236052 394670
rect 236000 394606 236052 394612
rect 236092 394052 236144 394058
rect 236092 393994 236144 394000
rect 236000 393984 236052 393990
rect 236000 393926 236052 393932
rect 235724 393848 235776 393854
rect 235724 393790 235776 393796
rect 235448 393712 235500 393718
rect 235448 393654 235500 393660
rect 235356 352708 235408 352714
rect 235356 352650 235408 352656
rect 235264 87780 235316 87786
rect 235264 87722 235316 87728
rect 235172 25696 235224 25702
rect 235172 25638 235224 25644
rect 235080 20324 235132 20330
rect 235080 20266 235132 20272
rect 234988 20256 235040 20262
rect 234988 20198 235040 20204
rect 234896 18692 234948 18698
rect 234896 18634 234948 18640
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 234620 6724 234672 6730
rect 234620 6666 234672 6672
rect 234894 5536 234950 5545
rect 234894 5471 234950 5480
rect 234908 4078 234936 5471
rect 234896 4072 234948 4078
rect 234896 4014 234948 4020
rect 235816 3936 235868 3942
rect 235816 3878 235868 3884
rect 234252 3732 234304 3738
rect 234252 3674 234304 3680
rect 234620 3120 234672 3126
rect 234620 3062 234672 3068
rect 234632 480 234660 3062
rect 235828 480 235856 3878
rect 236012 3777 236040 393926
rect 236104 3942 236132 393994
rect 236196 393922 236224 400044
rect 236288 394398 236316 400044
rect 236276 394392 236328 394398
rect 236276 394334 236328 394340
rect 236380 394058 236408 400044
rect 236368 394052 236420 394058
rect 236368 393994 236420 394000
rect 236184 393916 236236 393922
rect 236184 393858 236236 393864
rect 236472 393836 236500 400044
rect 236288 393808 236500 393836
rect 236288 393802 236316 393808
rect 236196 393774 236316 393802
rect 236196 6594 236224 393774
rect 236276 393712 236328 393718
rect 236276 393654 236328 393660
rect 236368 393712 236420 393718
rect 236368 393654 236420 393660
rect 236288 6662 236316 393654
rect 236276 6656 236328 6662
rect 236276 6598 236328 6604
rect 236184 6588 236236 6594
rect 236184 6530 236236 6536
rect 236380 6526 236408 393654
rect 236564 389174 236592 400044
rect 236656 393990 236684 400044
rect 236748 398177 236776 400044
rect 236734 398168 236790 398177
rect 236734 398103 236790 398112
rect 236736 394188 236788 394194
rect 236736 394130 236788 394136
rect 236644 393984 236696 393990
rect 236644 393926 236696 393932
rect 236748 389174 236776 394130
rect 236840 393786 236868 400044
rect 236828 393780 236880 393786
rect 236828 393722 236880 393728
rect 236932 393718 236960 400044
rect 237024 397186 237052 400044
rect 237116 397769 237144 400044
rect 237102 397760 237158 397769
rect 237102 397695 237158 397704
rect 237208 397497 237236 400044
rect 237300 397633 237328 400044
rect 237392 398002 237420 400044
rect 237380 397996 237432 398002
rect 237380 397938 237432 397944
rect 237286 397624 237342 397633
rect 237286 397559 237342 397568
rect 237194 397488 237250 397497
rect 237194 397423 237250 397432
rect 237012 397180 237064 397186
rect 237012 397122 237064 397128
rect 237380 394596 237432 394602
rect 237380 394538 237432 394544
rect 237392 393938 237420 394538
rect 237484 394040 237512 400044
rect 237576 394108 237604 400044
rect 237668 394505 237696 400044
rect 237654 394496 237710 394505
rect 237654 394431 237710 394440
rect 237760 394262 237788 400044
rect 237852 394641 237880 400044
rect 237944 394738 237972 400044
rect 237932 394732 237984 394738
rect 237932 394674 237984 394680
rect 237838 394632 237894 394641
rect 238036 394602 238064 400044
rect 237838 394567 237894 394576
rect 238024 394596 238076 394602
rect 238024 394538 238076 394544
rect 238022 394496 238078 394505
rect 238022 394431 238078 394440
rect 237748 394256 237800 394262
rect 237748 394198 237800 394204
rect 237576 394080 237788 394108
rect 237484 394012 237696 394040
rect 237392 393910 237512 393938
rect 237380 393848 237432 393854
rect 237380 393790 237432 393796
rect 236920 393712 236972 393718
rect 236920 393654 236972 393660
rect 236472 389146 236592 389174
rect 236656 389146 236776 389174
rect 236472 25634 236500 389146
rect 236460 25628 236512 25634
rect 236460 25570 236512 25576
rect 236368 6520 236420 6526
rect 236368 6462 236420 6468
rect 236092 3936 236144 3942
rect 236092 3878 236144 3884
rect 235998 3768 236054 3777
rect 235998 3703 236054 3712
rect 236552 3528 236604 3534
rect 236552 3470 236604 3476
rect 236564 3330 236592 3470
rect 236552 3324 236604 3330
rect 236552 3266 236604 3272
rect 236656 3194 236684 389146
rect 237392 9110 237420 393790
rect 237484 9178 237512 393910
rect 237564 393916 237616 393922
rect 237564 393858 237616 393864
rect 237576 9246 237604 393858
rect 237668 9314 237696 394012
rect 237760 20194 237788 394080
rect 237930 393952 237986 393961
rect 237930 393887 237986 393896
rect 237840 391264 237892 391270
rect 237840 391206 237892 391212
rect 237852 27198 237880 391206
rect 237944 27266 237972 393887
rect 238036 177478 238064 394431
rect 238128 351286 238156 400044
rect 238220 398138 238248 400044
rect 238208 398132 238260 398138
rect 238208 398074 238260 398080
rect 238208 397520 238260 397526
rect 238208 397462 238260 397468
rect 238220 391610 238248 397462
rect 238312 393854 238340 400044
rect 238404 397769 238432 400044
rect 238390 397760 238446 397769
rect 238390 397695 238446 397704
rect 238496 397633 238524 400044
rect 238482 397624 238538 397633
rect 238482 397559 238538 397568
rect 238588 397497 238616 400044
rect 238574 397488 238630 397497
rect 238574 397423 238630 397432
rect 238680 397089 238708 400044
rect 238772 397526 238800 400044
rect 238760 397520 238812 397526
rect 238760 397462 238812 397468
rect 238666 397080 238722 397089
rect 238666 397015 238722 397024
rect 238864 395214 238892 400044
rect 238852 395208 238904 395214
rect 238852 395150 238904 395156
rect 238392 394732 238444 394738
rect 238392 394674 238444 394680
rect 238300 393848 238352 393854
rect 238300 393790 238352 393796
rect 238208 391604 238260 391610
rect 238208 391546 238260 391552
rect 238404 391270 238432 394674
rect 238760 394460 238812 394466
rect 238760 394402 238812 394408
rect 238392 391264 238444 391270
rect 238392 391206 238444 391212
rect 238116 351280 238168 351286
rect 238116 351222 238168 351228
rect 238024 177472 238076 177478
rect 238024 177414 238076 177420
rect 238024 177336 238076 177342
rect 238024 177278 238076 177284
rect 237932 27260 237984 27266
rect 237932 27202 237984 27208
rect 237840 27192 237892 27198
rect 237840 27134 237892 27140
rect 237748 20188 237800 20194
rect 237748 20130 237800 20136
rect 238036 16574 238064 177278
rect 238036 16546 238156 16574
rect 237656 9308 237708 9314
rect 237656 9250 237708 9256
rect 237564 9240 237616 9246
rect 237564 9182 237616 9188
rect 237472 9172 237524 9178
rect 237472 9114 237524 9120
rect 237380 9104 237432 9110
rect 237380 9046 237432 9052
rect 237012 3664 237064 3670
rect 237012 3606 237064 3612
rect 236644 3188 236696 3194
rect 236644 3130 236696 3136
rect 237024 480 237052 3606
rect 238128 480 238156 16546
rect 238772 9042 238800 394402
rect 238852 394188 238904 394194
rect 238852 394130 238904 394136
rect 238864 10674 238892 394130
rect 238956 394108 238984 400044
rect 239048 394176 239076 400044
rect 239140 394466 239168 400044
rect 239232 394505 239260 400044
rect 239324 397662 239352 400044
rect 239312 397656 239364 397662
rect 239312 397598 239364 397604
rect 239218 394496 239274 394505
rect 239128 394460 239180 394466
rect 239218 394431 239274 394440
rect 239128 394402 239180 394408
rect 239416 394194 239444 400044
rect 239404 394188 239456 394194
rect 239048 394148 239260 394176
rect 238956 394080 239168 394108
rect 239034 393952 239090 393961
rect 239034 393887 239090 393896
rect 238944 392148 238996 392154
rect 238944 392090 238996 392096
rect 238852 10668 238904 10674
rect 238852 10610 238904 10616
rect 238956 10470 238984 392090
rect 239048 20058 239076 393887
rect 239140 20126 239168 394080
rect 239232 394040 239260 394148
rect 239404 394130 239456 394136
rect 239232 394012 239352 394040
rect 239220 390652 239272 390658
rect 239220 390594 239272 390600
rect 239128 20120 239180 20126
rect 239128 20062 239180 20068
rect 239036 20052 239088 20058
rect 239036 19994 239088 20000
rect 239232 19990 239260 390594
rect 239324 27130 239352 394012
rect 239508 390658 239536 400044
rect 239496 390652 239548 390658
rect 239496 390594 239548 390600
rect 239600 389174 239628 400044
rect 239692 392154 239720 400044
rect 239784 397497 239812 400044
rect 239876 397934 239904 400044
rect 239864 397928 239916 397934
rect 239864 397870 239916 397876
rect 239864 397792 239916 397798
rect 239864 397734 239916 397740
rect 239770 397488 239826 397497
rect 239770 397423 239826 397432
rect 239772 395208 239824 395214
rect 239772 395150 239824 395156
rect 239680 392148 239732 392154
rect 239680 392090 239732 392096
rect 239784 391542 239812 395150
rect 239876 392834 239904 397734
rect 239968 397497 239996 400044
rect 240060 397633 240088 400044
rect 240046 397624 240102 397633
rect 240046 397559 240102 397568
rect 239954 397488 240010 397497
rect 239954 397423 240010 397432
rect 240152 394330 240180 400044
rect 240244 397798 240272 400044
rect 240232 397792 240284 397798
rect 240232 397734 240284 397740
rect 240140 394324 240192 394330
rect 240140 394266 240192 394272
rect 240140 394188 240192 394194
rect 240140 394130 240192 394136
rect 239864 392828 239916 392834
rect 239864 392770 239916 392776
rect 239772 391536 239824 391542
rect 239772 391478 239824 391484
rect 239416 389146 239628 389174
rect 239416 87718 239444 389146
rect 239404 87712 239456 87718
rect 239404 87654 239456 87660
rect 239312 27124 239364 27130
rect 239312 27066 239364 27072
rect 239220 19984 239272 19990
rect 239220 19926 239272 19932
rect 240152 12170 240180 394130
rect 240232 394120 240284 394126
rect 240232 394062 240284 394068
rect 240244 17474 240272 394062
rect 240336 394058 240364 400044
rect 240324 394052 240376 394058
rect 240428 394040 240456 400044
rect 240520 397866 240548 400044
rect 240508 397860 240560 397866
rect 240508 397802 240560 397808
rect 240612 394126 240640 400044
rect 240704 394194 240732 400044
rect 240796 399945 240824 400044
rect 240782 399936 240838 399945
rect 240782 399871 240838 399880
rect 240692 394188 240744 394194
rect 240692 394130 240744 394136
rect 240600 394120 240652 394126
rect 240600 394062 240652 394068
rect 240692 394052 240744 394058
rect 240428 394012 240548 394040
rect 240324 393994 240376 394000
rect 240416 393916 240468 393922
rect 240416 393858 240468 393864
rect 240324 393848 240376 393854
rect 240324 393790 240376 393796
rect 240336 21690 240364 393790
rect 240428 26994 240456 393858
rect 240520 27062 240548 394012
rect 240692 393994 240744 394000
rect 240600 393984 240652 393990
rect 240600 393926 240652 393932
rect 240612 177410 240640 393926
rect 240704 352646 240732 393994
rect 240888 389910 240916 400044
rect 240876 389904 240928 389910
rect 240876 389846 240928 389852
rect 240980 389174 241008 400044
rect 241072 393990 241100 400044
rect 241060 393984 241112 393990
rect 241060 393926 241112 393932
rect 241164 393854 241192 400044
rect 241256 393922 241284 400044
rect 241348 397497 241376 400044
rect 241334 397488 241390 397497
rect 241334 397423 241390 397432
rect 241440 396953 241468 400044
rect 241532 398206 241560 400044
rect 241520 398200 241572 398206
rect 241520 398142 241572 398148
rect 241520 398064 241572 398070
rect 241520 398006 241572 398012
rect 241426 396944 241482 396953
rect 241426 396879 241482 396888
rect 241532 395622 241560 398006
rect 241624 395894 241652 400044
rect 241716 397050 241744 400044
rect 241704 397044 241756 397050
rect 241704 396986 241756 396992
rect 241808 396074 241836 400044
rect 241716 396046 241836 396074
rect 241612 395888 241664 395894
rect 241612 395830 241664 395836
rect 241520 395616 241572 395622
rect 241520 395558 241572 395564
rect 241520 394120 241572 394126
rect 241520 394062 241572 394068
rect 241244 393916 241296 393922
rect 241244 393858 241296 393864
rect 241152 393848 241204 393854
rect 241152 393790 241204 393796
rect 240888 389146 241008 389174
rect 240888 354210 240916 389146
rect 240876 354204 240928 354210
rect 240876 354146 240928 354152
rect 240784 354068 240836 354074
rect 240784 354010 240836 354016
rect 240692 352640 240744 352646
rect 240692 352582 240744 352588
rect 240600 177404 240652 177410
rect 240600 177346 240652 177352
rect 240508 27056 240560 27062
rect 240508 26998 240560 27004
rect 240416 26988 240468 26994
rect 240416 26930 240468 26936
rect 240324 21684 240376 21690
rect 240324 21626 240376 21632
rect 240232 17468 240284 17474
rect 240232 17410 240284 17416
rect 240140 12164 240192 12170
rect 240140 12106 240192 12112
rect 238944 10464 238996 10470
rect 238944 10406 238996 10412
rect 238760 9036 238812 9042
rect 238760 8978 238812 8984
rect 239404 4140 239456 4146
rect 239404 4082 239456 4088
rect 239416 3942 239444 4082
rect 239312 3936 239364 3942
rect 239312 3878 239364 3884
rect 239404 3936 239456 3942
rect 239404 3878 239456 3884
rect 239324 3754 239352 3878
rect 239324 3726 239536 3754
rect 239508 3670 239536 3726
rect 239496 3664 239548 3670
rect 239310 3632 239366 3641
rect 239496 3606 239548 3612
rect 239310 3567 239366 3576
rect 239324 480 239352 3567
rect 239404 3528 239456 3534
rect 239404 3470 239456 3476
rect 240506 3496 240562 3505
rect 239416 3330 239444 3470
rect 240506 3431 240562 3440
rect 239404 3324 239456 3330
rect 239404 3266 239456 3272
rect 240520 480 240548 3431
rect 240796 3330 240824 354010
rect 241532 10402 241560 394062
rect 241612 393984 241664 393990
rect 241612 393926 241664 393932
rect 241716 393938 241744 396046
rect 241900 394126 241928 400044
rect 241888 394120 241940 394126
rect 241888 394062 241940 394068
rect 241520 10396 241572 10402
rect 241520 10338 241572 10344
rect 241624 10334 241652 393926
rect 241716 393910 241836 393938
rect 241704 393848 241756 393854
rect 241704 393790 241756 393796
rect 241716 21622 241744 393790
rect 241808 26926 241836 393910
rect 241888 393916 241940 393922
rect 241888 393858 241940 393864
rect 241900 87650 241928 393858
rect 241992 393854 242020 400044
rect 242084 397594 242112 400044
rect 242072 397588 242124 397594
rect 242072 397530 242124 397536
rect 242072 397112 242124 397118
rect 242072 397054 242124 397060
rect 241980 393848 242032 393854
rect 241980 393790 242032 393796
rect 242084 389174 242112 397054
rect 242176 393990 242204 400044
rect 242268 396846 242296 400044
rect 242256 396840 242308 396846
rect 242256 396782 242308 396788
rect 242164 393984 242216 393990
rect 242164 393926 242216 393932
rect 242360 393922 242388 400044
rect 242452 397633 242480 400044
rect 242544 397769 242572 400044
rect 242636 398818 242664 400044
rect 242624 398812 242676 398818
rect 242624 398754 242676 398760
rect 242624 397928 242676 397934
rect 242624 397870 242676 397876
rect 242530 397760 242586 397769
rect 242530 397695 242586 397704
rect 242438 397624 242494 397633
rect 242438 397559 242494 397568
rect 242440 395888 242492 395894
rect 242440 395830 242492 395836
rect 242348 393916 242400 393922
rect 242348 393858 242400 393864
rect 242452 392698 242480 395830
rect 242440 392692 242492 392698
rect 242440 392634 242492 392640
rect 242636 389174 242664 397870
rect 242728 397497 242756 400044
rect 242820 397905 242848 400044
rect 242806 397896 242862 397905
rect 242806 397831 242862 397840
rect 242714 397488 242770 397497
rect 242714 397423 242770 397432
rect 242084 389146 242204 389174
rect 241888 87644 241940 87650
rect 241888 87586 241940 87592
rect 241796 26920 241848 26926
rect 241796 26862 241848 26868
rect 241704 21616 241756 21622
rect 241704 21558 241756 21564
rect 241612 10328 241664 10334
rect 241612 10270 241664 10276
rect 241704 4956 241756 4962
rect 241704 4898 241756 4904
rect 240784 3324 240836 3330
rect 240784 3266 240836 3272
rect 241716 480 241744 4898
rect 242176 4146 242204 389146
rect 242452 389146 242664 389174
rect 242452 10538 242480 389146
rect 242440 10532 242492 10538
rect 242440 10474 242492 10480
rect 242912 6458 242940 400044
rect 242900 6452 242952 6458
rect 242900 6394 242952 6400
rect 243004 6390 243032 400044
rect 243096 393922 243124 400044
rect 243188 397730 243216 400044
rect 243176 397724 243228 397730
rect 243176 397666 243228 397672
rect 243176 394256 243228 394262
rect 243176 394198 243228 394204
rect 243084 393916 243136 393922
rect 243084 393858 243136 393864
rect 243188 393802 243216 394198
rect 243096 393774 243216 393802
rect 243096 12034 243124 393774
rect 243176 393712 243228 393718
rect 243176 393654 243228 393660
rect 243084 12028 243136 12034
rect 243084 11970 243136 11976
rect 243188 11966 243216 393654
rect 243280 12102 243308 400044
rect 243372 394194 243400 400044
rect 243360 394188 243412 394194
rect 243360 394130 243412 394136
rect 243464 394040 243492 400044
rect 243556 394262 243584 400044
rect 243544 394256 243596 394262
rect 243544 394198 243596 394204
rect 243648 394040 243676 400044
rect 243740 398070 243768 400044
rect 243728 398064 243780 398070
rect 243728 398006 243780 398012
rect 243728 394188 243780 394194
rect 243728 394130 243780 394136
rect 243372 394012 243492 394040
rect 243556 394012 243676 394040
rect 243372 13530 243400 394012
rect 243452 393916 243504 393922
rect 243452 393858 243504 393864
rect 243464 82210 243492 393858
rect 243556 86562 243584 394012
rect 243740 389174 243768 394130
rect 243832 393718 243860 400044
rect 243924 398993 243952 400044
rect 243910 398984 243966 398993
rect 243910 398919 243966 398928
rect 243912 397996 243964 398002
rect 243912 397938 243964 397944
rect 243924 394262 243952 397938
rect 244016 397497 244044 400044
rect 244108 397633 244136 400044
rect 244200 397769 244228 400044
rect 244292 397934 244320 400044
rect 244384 399022 244412 400044
rect 244372 399016 244424 399022
rect 244372 398958 244424 398964
rect 244370 398712 244426 398721
rect 244370 398647 244426 398656
rect 244280 397928 244332 397934
rect 244280 397870 244332 397876
rect 244186 397760 244242 397769
rect 244186 397695 244242 397704
rect 244094 397624 244150 397633
rect 244094 397559 244150 397568
rect 244002 397488 244058 397497
rect 244002 397423 244058 397432
rect 244384 396817 244412 398647
rect 244370 396808 244426 396817
rect 244370 396743 244426 396752
rect 244004 394664 244056 394670
rect 244004 394606 244056 394612
rect 244016 394398 244044 394606
rect 244004 394392 244056 394398
rect 244004 394334 244056 394340
rect 243912 394256 243964 394262
rect 243912 394198 243964 394204
rect 244372 394188 244424 394194
rect 244372 394130 244424 394136
rect 244280 394120 244332 394126
rect 244280 394062 244332 394068
rect 244186 393816 244242 393825
rect 244186 393751 244188 393760
rect 244240 393751 244242 393760
rect 244188 393722 244240 393728
rect 243820 393712 243872 393718
rect 243820 393654 243872 393660
rect 243648 389146 243768 389174
rect 243648 352578 243676 389146
rect 243636 352572 243688 352578
rect 243636 352514 243688 352520
rect 243544 86556 243596 86562
rect 243544 86498 243596 86504
rect 243452 82204 243504 82210
rect 243452 82146 243504 82152
rect 243360 13524 243412 13530
rect 243360 13466 243412 13472
rect 243268 12096 243320 12102
rect 243268 12038 243320 12044
rect 243176 11960 243228 11966
rect 243176 11902 243228 11908
rect 244292 11898 244320 394062
rect 244280 11892 244332 11898
rect 244280 11834 244332 11840
rect 244384 11830 244412 394130
rect 244476 393938 244504 400044
rect 244568 394040 244596 400044
rect 244660 395146 244688 400044
rect 244648 395140 244700 395146
rect 244648 395082 244700 395088
rect 244648 394052 244700 394058
rect 244568 394012 244648 394040
rect 244648 393994 244700 394000
rect 244476 393910 244688 393938
rect 244464 393848 244516 393854
rect 244464 393790 244516 393796
rect 244476 21486 244504 393790
rect 244556 393780 244608 393786
rect 244556 393722 244608 393728
rect 244464 21480 244516 21486
rect 244464 21422 244516 21428
rect 244568 21418 244596 393722
rect 244660 21554 244688 393910
rect 244752 393854 244780 400044
rect 244844 398954 244872 400044
rect 244832 398948 244884 398954
rect 244832 398890 244884 398896
rect 244832 397520 244884 397526
rect 244832 397462 244884 397468
rect 244740 393848 244792 393854
rect 244740 393790 244792 393796
rect 244740 393712 244792 393718
rect 244740 393654 244792 393660
rect 244752 355434 244780 393654
rect 244844 393650 244872 397462
rect 244936 394126 244964 400044
rect 244924 394120 244976 394126
rect 244924 394062 244976 394068
rect 245028 393718 245056 400044
rect 245016 393712 245068 393718
rect 245016 393654 245068 393660
rect 244832 393644 244884 393650
rect 244832 393586 244884 393592
rect 245120 393530 245148 400044
rect 245212 394194 245240 400044
rect 245200 394188 245252 394194
rect 245200 394130 245252 394136
rect 245200 394052 245252 394058
rect 245200 393994 245252 394000
rect 244844 393502 245148 393530
rect 244740 355428 244792 355434
rect 244740 355370 244792 355376
rect 244740 354000 244792 354006
rect 244740 353942 244792 353948
rect 244648 21548 244700 21554
rect 244648 21490 244700 21496
rect 244556 21412 244608 21418
rect 244556 21354 244608 21360
rect 244752 16574 244780 353942
rect 244844 86494 244872 393502
rect 244924 393440 244976 393446
rect 244924 393382 244976 393388
rect 244832 86488 244884 86494
rect 244832 86430 244884 86436
rect 244936 82278 244964 393382
rect 245212 386414 245240 393994
rect 245304 393786 245332 400044
rect 245396 398002 245424 400044
rect 245384 397996 245436 398002
rect 245384 397938 245436 397944
rect 245488 397497 245516 400044
rect 245474 397488 245530 397497
rect 245474 397423 245530 397432
rect 245580 396681 245608 400044
rect 245566 396672 245622 396681
rect 245566 396607 245622 396616
rect 245384 395140 245436 395146
rect 245384 395082 245436 395088
rect 245292 393780 245344 393786
rect 245292 393722 245344 393728
rect 245396 391406 245424 395082
rect 245672 392426 245700 400044
rect 245660 392420 245712 392426
rect 245660 392362 245712 392368
rect 245764 392306 245792 400044
rect 245672 392278 245792 392306
rect 245384 391400 245436 391406
rect 245384 391342 245436 391348
rect 245028 386386 245240 386414
rect 245028 354142 245056 386386
rect 245016 354136 245068 354142
rect 245016 354078 245068 354084
rect 244924 82272 244976 82278
rect 244924 82214 244976 82220
rect 244752 16546 245240 16574
rect 244372 11824 244424 11830
rect 244372 11766 244424 11772
rect 242992 6384 243044 6390
rect 242992 6326 243044 6332
rect 242164 4140 242216 4146
rect 242164 4082 242216 4088
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242900 3188 242952 3194
rect 242900 3130 242952 3136
rect 242912 480 242940 3130
rect 244108 480 244136 3334
rect 245212 480 245240 16546
rect 245672 11762 245700 392278
rect 245752 392216 245804 392222
rect 245752 392158 245804 392164
rect 245764 13394 245792 392158
rect 245856 391338 245884 400044
rect 245948 398886 245976 400044
rect 245936 398880 245988 398886
rect 245936 398822 245988 398828
rect 246040 392170 246068 400044
rect 245948 392142 246068 392170
rect 245844 391332 245896 391338
rect 245844 391274 245896 391280
rect 245844 391060 245896 391066
rect 245844 391002 245896 391008
rect 245752 13388 245804 13394
rect 245752 13330 245804 13336
rect 245856 13326 245884 391002
rect 245948 13462 245976 392142
rect 246132 392034 246160 400044
rect 246224 398546 246252 400044
rect 246212 398540 246264 398546
rect 246212 398482 246264 398488
rect 246212 394188 246264 394194
rect 246212 394130 246264 394136
rect 246224 393825 246252 394130
rect 246210 393816 246266 393825
rect 246210 393751 246266 393760
rect 246212 392420 246264 392426
rect 246212 392362 246264 392368
rect 246040 392006 246160 392034
rect 246040 23186 246068 392006
rect 246120 390108 246172 390114
rect 246120 390050 246172 390056
rect 246028 23180 246080 23186
rect 246028 23122 246080 23128
rect 246132 23118 246160 390050
rect 246224 86426 246252 392362
rect 246316 392222 246344 400044
rect 246304 392216 246356 392222
rect 246304 392158 246356 392164
rect 246408 390114 246436 400044
rect 246500 398313 246528 400044
rect 246486 398304 246542 398313
rect 246486 398239 246542 398248
rect 246488 398132 246540 398138
rect 246488 398074 246540 398080
rect 246396 390108 246448 390114
rect 246396 390050 246448 390056
rect 246500 389174 246528 398074
rect 246592 391066 246620 400044
rect 246684 397633 246712 400044
rect 246776 398478 246804 400044
rect 246764 398472 246816 398478
rect 246764 398414 246816 398420
rect 246670 397624 246726 397633
rect 246670 397559 246726 397568
rect 246868 397497 246896 400044
rect 246960 397769 246988 400044
rect 246946 397760 247002 397769
rect 246946 397695 247002 397704
rect 246948 397656 247000 397662
rect 246948 397598 247000 397604
rect 246854 397488 246910 397497
rect 246854 397423 246910 397432
rect 246960 394126 246988 397598
rect 246948 394120 247000 394126
rect 246948 394062 247000 394068
rect 247052 393854 247080 400044
rect 247040 393848 247092 393854
rect 247040 393790 247092 393796
rect 247144 392170 247172 400044
rect 247236 396778 247264 400044
rect 247328 398342 247356 400044
rect 247316 398336 247368 398342
rect 247316 398278 247368 398284
rect 247316 397928 247368 397934
rect 247316 397870 247368 397876
rect 247328 397662 247356 397870
rect 247316 397656 247368 397662
rect 247316 397598 247368 397604
rect 247224 396772 247276 396778
rect 247224 396714 247276 396720
rect 247420 393938 247448 400044
rect 247052 392142 247172 392170
rect 247236 393910 247448 393938
rect 246580 391060 246632 391066
rect 246580 391002 246632 391008
rect 246500 389146 246620 389174
rect 246592 354278 246620 389146
rect 246580 354272 246632 354278
rect 246580 354214 246632 354220
rect 246212 86420 246264 86426
rect 246212 86362 246264 86368
rect 246120 23112 246172 23118
rect 246120 23054 246172 23060
rect 245936 13456 245988 13462
rect 245936 13398 245988 13404
rect 245844 13320 245896 13326
rect 245844 13262 245896 13268
rect 247052 13258 247080 392142
rect 247132 392080 247184 392086
rect 247132 392022 247184 392028
rect 247040 13252 247092 13258
rect 247040 13194 247092 13200
rect 247144 13122 247172 392022
rect 247236 13190 247264 393910
rect 247316 393848 247368 393854
rect 247316 393790 247368 393796
rect 247408 393848 247460 393854
rect 247408 393790 247460 393796
rect 247328 18630 247356 393790
rect 247420 22982 247448 393790
rect 247512 23050 247540 400044
rect 247604 86358 247632 400044
rect 247696 398138 247724 400044
rect 247684 398132 247736 398138
rect 247684 398074 247736 398080
rect 247684 397792 247736 397798
rect 247684 397734 247736 397740
rect 247592 86352 247644 86358
rect 247592 86294 247644 86300
rect 247500 23044 247552 23050
rect 247500 22986 247552 22992
rect 247408 22976 247460 22982
rect 247408 22918 247460 22924
rect 247316 18624 247368 18630
rect 247316 18566 247368 18572
rect 247224 13184 247276 13190
rect 247224 13126 247276 13132
rect 247132 13116 247184 13122
rect 247132 13058 247184 13064
rect 245660 11756 245712 11762
rect 245660 11698 245712 11704
rect 247696 10606 247724 397734
rect 247788 392086 247816 400044
rect 247880 393854 247908 400044
rect 247972 398041 248000 400044
rect 247958 398032 248014 398041
rect 247958 397967 248014 397976
rect 247960 397860 248012 397866
rect 247960 397802 248012 397808
rect 247868 393848 247920 393854
rect 247868 393790 247920 393796
rect 247776 392080 247828 392086
rect 247776 392022 247828 392028
rect 247972 391474 248000 397802
rect 248064 397633 248092 400044
rect 248156 397769 248184 400044
rect 248142 397760 248198 397769
rect 248142 397695 248198 397704
rect 248050 397624 248106 397633
rect 248050 397559 248106 397568
rect 248248 397497 248276 400044
rect 248340 397905 248368 400044
rect 248326 397896 248382 397905
rect 248326 397831 248382 397840
rect 248234 397488 248290 397497
rect 248234 397423 248290 397432
rect 248432 392086 248460 400044
rect 248524 399129 248552 400044
rect 248510 399120 248566 399129
rect 248510 399055 248566 399064
rect 248512 398200 248564 398206
rect 248512 398142 248564 398148
rect 248524 397866 248552 398142
rect 248512 397860 248564 397866
rect 248512 397802 248564 397808
rect 248512 395888 248564 395894
rect 248512 395830 248564 395836
rect 248420 392080 248472 392086
rect 248420 392022 248472 392028
rect 248420 391944 248472 391950
rect 248420 391886 248472 391892
rect 247960 391468 248012 391474
rect 247960 391410 248012 391416
rect 247684 10600 247736 10606
rect 247684 10542 247736 10548
rect 246396 3596 246448 3602
rect 246396 3538 246448 3544
rect 246408 480 246436 3538
rect 248432 3534 248460 391886
rect 248524 14754 248552 395830
rect 248616 14890 248644 400044
rect 248708 393854 248736 400044
rect 248800 398585 248828 400044
rect 248786 398576 248842 398585
rect 248786 398511 248842 398520
rect 248696 393848 248748 393854
rect 248696 393790 248748 393796
rect 248892 392170 248920 400044
rect 248984 393938 249012 400044
rect 249076 395706 249104 400044
rect 249168 395894 249196 400044
rect 249260 395894 249288 400044
rect 249156 395888 249208 395894
rect 249156 395830 249208 395836
rect 249248 395888 249300 395894
rect 249248 395830 249300 395836
rect 249076 395678 249288 395706
rect 248984 393910 249104 393938
rect 248972 393848 249024 393854
rect 248972 393790 249024 393796
rect 248800 392142 248920 392170
rect 248696 392012 248748 392018
rect 248696 391954 248748 391960
rect 248604 14884 248656 14890
rect 248604 14826 248656 14832
rect 248512 14748 248564 14754
rect 248512 14690 248564 14696
rect 248708 14686 248736 391954
rect 248800 14822 248828 392142
rect 248880 392080 248932 392086
rect 248880 392022 248932 392028
rect 248892 22914 248920 392022
rect 248880 22908 248932 22914
rect 248880 22850 248932 22856
rect 248984 22846 249012 393790
rect 249076 177342 249104 393910
rect 249260 392630 249288 395678
rect 249248 392624 249300 392630
rect 249248 392566 249300 392572
rect 249352 391950 249380 400044
rect 249444 392018 249472 400044
rect 249536 397633 249564 400044
rect 249522 397624 249578 397633
rect 249522 397559 249578 397568
rect 249628 397497 249656 400044
rect 249720 397769 249748 400044
rect 249706 397760 249762 397769
rect 249706 397695 249762 397704
rect 249614 397488 249670 397497
rect 249614 397423 249670 397432
rect 249524 395888 249576 395894
rect 249524 395830 249576 395836
rect 249432 392012 249484 392018
rect 249432 391954 249484 391960
rect 249340 391944 249392 391950
rect 249340 391886 249392 391892
rect 249536 389842 249564 395830
rect 249812 392086 249840 400044
rect 249904 398177 249932 400044
rect 249890 398168 249946 398177
rect 249890 398103 249946 398112
rect 249892 394052 249944 394058
rect 249892 393994 249944 394000
rect 249800 392080 249852 392086
rect 249800 392022 249852 392028
rect 249800 391944 249852 391950
rect 249800 391886 249852 391892
rect 249524 389836 249576 389842
rect 249524 389778 249576 389784
rect 249064 177336 249116 177342
rect 249064 177278 249116 177284
rect 248972 22840 249024 22846
rect 248972 22782 249024 22788
rect 248788 14816 248840 14822
rect 248788 14758 248840 14764
rect 248696 14680 248748 14686
rect 248696 14622 248748 14628
rect 249812 5234 249840 391886
rect 249904 14482 249932 393994
rect 249996 393938 250024 400044
rect 250088 394074 250116 400044
rect 250180 398857 250208 400044
rect 250166 398848 250222 398857
rect 250166 398783 250222 398792
rect 250168 398744 250220 398750
rect 250168 398686 250220 398692
rect 250180 397866 250208 398686
rect 250168 397860 250220 397866
rect 250168 397802 250220 397808
rect 250088 394046 250208 394074
rect 249996 393910 250116 393938
rect 249984 393848 250036 393854
rect 249984 393790 250036 393796
rect 249996 14550 250024 393790
rect 250088 14618 250116 393910
rect 250180 393394 250208 394046
rect 250272 393854 250300 400044
rect 250260 393848 250312 393854
rect 250260 393790 250312 393796
rect 250364 393666 250392 400044
rect 250456 393938 250484 400044
rect 250548 394058 250576 400044
rect 250536 394052 250588 394058
rect 250536 393994 250588 394000
rect 250456 393910 250576 393938
rect 250364 393638 250484 393666
rect 250180 393366 250392 393394
rect 250260 392148 250312 392154
rect 250260 392090 250312 392096
rect 250168 392080 250220 392086
rect 250168 392022 250220 392028
rect 250180 22778 250208 392022
rect 250272 24410 250300 392090
rect 250364 24478 250392 393366
rect 250456 392154 250484 393638
rect 250444 392148 250496 392154
rect 250444 392090 250496 392096
rect 250444 389360 250496 389366
rect 250444 389302 250496 389308
rect 250456 86290 250484 389302
rect 250548 355366 250576 393910
rect 250640 389366 250668 400044
rect 250732 391950 250760 400044
rect 250824 397633 250852 400044
rect 250916 397905 250944 400044
rect 250902 397896 250958 397905
rect 250902 397831 250958 397840
rect 250810 397624 250866 397633
rect 250810 397559 250866 397568
rect 251008 397497 251036 400044
rect 251100 397769 251128 400044
rect 251086 397760 251142 397769
rect 251086 397695 251142 397704
rect 250810 397488 250866 397497
rect 250810 397423 250866 397432
rect 250994 397488 251050 397497
rect 250994 397423 251050 397432
rect 250720 391944 250772 391950
rect 250720 391886 250772 391892
rect 250824 391270 250852 397423
rect 251192 393854 251220 400044
rect 251284 398313 251312 400044
rect 251270 398304 251326 398313
rect 251270 398239 251326 398248
rect 251272 394596 251324 394602
rect 251272 394538 251324 394544
rect 251180 393848 251232 393854
rect 251180 393790 251232 393796
rect 251284 393802 251312 394538
rect 251376 393938 251404 400044
rect 251468 394074 251496 400044
rect 251560 397186 251588 400044
rect 251548 397180 251600 397186
rect 251548 397122 251600 397128
rect 251652 394602 251680 400044
rect 251640 394596 251692 394602
rect 251640 394538 251692 394544
rect 251468 394046 251680 394074
rect 251548 393984 251600 393990
rect 251376 393910 251496 393938
rect 251548 393926 251600 393932
rect 251284 393774 251404 393802
rect 251180 393712 251232 393718
rect 251180 393654 251232 393660
rect 250812 391264 250864 391270
rect 250812 391206 250864 391212
rect 250628 389360 250680 389366
rect 250628 389302 250680 389308
rect 250536 355360 250588 355366
rect 250536 355302 250588 355308
rect 250444 86284 250496 86290
rect 250444 86226 250496 86232
rect 250352 24472 250404 24478
rect 250352 24414 250404 24420
rect 250260 24404 250312 24410
rect 250260 24346 250312 24352
rect 250168 22772 250220 22778
rect 250168 22714 250220 22720
rect 250076 14612 250128 14618
rect 250076 14554 250128 14560
rect 249984 14544 250036 14550
rect 249984 14486 250036 14492
rect 249892 14476 249944 14482
rect 249892 14418 249944 14424
rect 249800 5228 249852 5234
rect 249800 5170 249852 5176
rect 251192 5166 251220 393654
rect 251272 390516 251324 390522
rect 251272 390458 251324 390464
rect 251180 5160 251232 5166
rect 251180 5102 251232 5108
rect 251284 5098 251312 390458
rect 251376 16114 251404 393774
rect 251468 16182 251496 393910
rect 251560 24206 251588 393926
rect 251652 24274 251680 394046
rect 251744 393990 251772 400044
rect 251732 393984 251784 393990
rect 251732 393926 251784 393932
rect 251732 393848 251784 393854
rect 251732 393790 251784 393796
rect 251744 24342 251772 393790
rect 251836 393718 251864 400044
rect 251824 393712 251876 393718
rect 251824 393654 251876 393660
rect 251928 389174 251956 400044
rect 252020 395554 252048 400044
rect 252008 395548 252060 395554
rect 252008 395490 252060 395496
rect 252112 390522 252140 400044
rect 252204 397905 252232 400044
rect 252190 397896 252246 397905
rect 252190 397831 252246 397840
rect 252296 397769 252324 400044
rect 252282 397760 252338 397769
rect 252282 397695 252338 397704
rect 252388 397497 252416 400044
rect 252480 397633 252508 400044
rect 252572 399265 252600 400044
rect 252664 399838 252692 400044
rect 252652 399832 252704 399838
rect 252652 399774 252704 399780
rect 252652 399696 252704 399702
rect 252652 399638 252704 399644
rect 252558 399256 252614 399265
rect 252558 399191 252614 399200
rect 252664 398970 252692 399638
rect 252572 398942 252692 398970
rect 252466 397624 252522 397633
rect 252466 397559 252522 397568
rect 252374 397488 252430 397497
rect 252374 397423 252430 397432
rect 252100 390516 252152 390522
rect 252100 390458 252152 390464
rect 251836 389146 251956 389174
rect 251836 354074 251864 389146
rect 251824 354068 251876 354074
rect 251824 354010 251876 354016
rect 251732 24336 251784 24342
rect 251732 24278 251784 24284
rect 251640 24268 251692 24274
rect 251640 24210 251692 24216
rect 251548 24200 251600 24206
rect 251548 24142 251600 24148
rect 251456 16176 251508 16182
rect 251456 16118 251508 16124
rect 251364 16108 251416 16114
rect 251364 16050 251416 16056
rect 251272 5092 251324 5098
rect 251272 5034 251324 5040
rect 252572 4962 252600 398942
rect 252650 398848 252706 398857
rect 252756 398818 252784 400044
rect 252650 398783 252706 398792
rect 252744 398812 252796 398818
rect 252664 395486 252692 398783
rect 252744 398754 252796 398760
rect 252742 398712 252798 398721
rect 252742 398647 252798 398656
rect 252652 395480 252704 395486
rect 252652 395422 252704 395428
rect 252652 393984 252704 393990
rect 252652 393926 252704 393932
rect 252664 5030 252692 393926
rect 252652 5024 252704 5030
rect 252652 4966 252704 4972
rect 252560 4956 252612 4962
rect 252560 4898 252612 4904
rect 252756 4894 252784 398647
rect 252848 394058 252876 400044
rect 252836 394052 252888 394058
rect 252836 393994 252888 394000
rect 252940 393990 252968 400044
rect 252928 393984 252980 393990
rect 252928 393926 252980 393932
rect 252928 393848 252980 393854
rect 252928 393790 252980 393796
rect 252836 393780 252888 393786
rect 252836 393722 252888 393728
rect 252848 7614 252876 393722
rect 252940 15910 252968 393790
rect 253032 15978 253060 400044
rect 253124 399430 253152 400044
rect 253216 399702 253244 400044
rect 253204 399696 253256 399702
rect 253204 399638 253256 399644
rect 253204 399560 253256 399566
rect 253204 399502 253256 399508
rect 253112 399424 253164 399430
rect 253112 399366 253164 399372
rect 253112 398812 253164 398818
rect 253112 398754 253164 398760
rect 253124 16046 253152 398754
rect 253216 397497 253244 399502
rect 253202 397488 253258 397497
rect 253202 397423 253258 397432
rect 253204 394052 253256 394058
rect 253204 393994 253256 394000
rect 253216 354006 253244 393994
rect 253308 393854 253336 400044
rect 253296 393848 253348 393854
rect 253296 393790 253348 393796
rect 253400 393786 253428 400044
rect 253492 399945 253520 400044
rect 253478 399936 253534 399945
rect 253478 399871 253534 399880
rect 253480 399832 253532 399838
rect 253480 399774 253532 399780
rect 253492 398954 253520 399774
rect 253480 398948 253532 398954
rect 253480 398890 253532 398896
rect 253480 398540 253532 398546
rect 253480 398482 253532 398488
rect 253492 398002 253520 398482
rect 253480 397996 253532 398002
rect 253480 397938 253532 397944
rect 253584 397497 253612 400044
rect 253676 399566 253704 400044
rect 253664 399560 253716 399566
rect 253664 399502 253716 399508
rect 253664 399424 253716 399430
rect 253664 399366 253716 399372
rect 253570 397488 253626 397497
rect 253570 397423 253626 397432
rect 253676 395418 253704 399366
rect 253768 397769 253796 400044
rect 253860 398449 253888 400044
rect 253846 398440 253902 398449
rect 253846 398375 253902 398384
rect 253754 397760 253810 397769
rect 253754 397695 253810 397704
rect 253952 396166 253980 400044
rect 254044 398041 254072 400044
rect 254030 398032 254086 398041
rect 254030 397967 254086 397976
rect 254032 396704 254084 396710
rect 254032 396646 254084 396652
rect 253940 396160 253992 396166
rect 253940 396102 253992 396108
rect 253664 395412 253716 395418
rect 253664 395354 253716 395360
rect 253388 393780 253440 393786
rect 253388 393722 253440 393728
rect 253204 354000 253256 354006
rect 253204 353942 253256 353948
rect 253112 16040 253164 16046
rect 253112 15982 253164 15988
rect 253020 15972 253072 15978
rect 253020 15914 253072 15920
rect 252928 15904 252980 15910
rect 252928 15846 252980 15852
rect 252836 7608 252888 7614
rect 252836 7550 252888 7556
rect 254044 6186 254072 396646
rect 254136 396574 254164 400044
rect 254228 397050 254256 400044
rect 254320 398886 254348 400044
rect 254308 398880 254360 398886
rect 254308 398822 254360 398828
rect 254216 397044 254268 397050
rect 254216 396986 254268 396992
rect 254412 396658 254440 400044
rect 254228 396630 254440 396658
rect 254124 396568 254176 396574
rect 254124 396510 254176 396516
rect 254124 396364 254176 396370
rect 254124 396306 254176 396312
rect 254136 6254 254164 396306
rect 254228 17338 254256 396630
rect 254400 396568 254452 396574
rect 254400 396510 254452 396516
rect 254308 396432 254360 396438
rect 254308 396374 254360 396380
rect 254216 17332 254268 17338
rect 254216 17274 254268 17280
rect 254320 17270 254348 396374
rect 254412 17406 254440 396510
rect 254504 24138 254532 400044
rect 254596 396370 254624 400044
rect 254688 396438 254716 400044
rect 254676 396432 254728 396438
rect 254676 396374 254728 396380
rect 254584 396364 254636 396370
rect 254584 396306 254636 396312
rect 254780 393990 254808 400044
rect 254872 396710 254900 400044
rect 254860 396704 254912 396710
rect 254860 396646 254912 396652
rect 254964 396250 254992 400044
rect 255056 397769 255084 400044
rect 255042 397760 255098 397769
rect 255042 397695 255098 397704
rect 255148 397633 255176 400044
rect 255240 397905 255268 400044
rect 255226 397896 255282 397905
rect 255226 397831 255282 397840
rect 255134 397624 255190 397633
rect 255134 397559 255190 397568
rect 255044 397044 255096 397050
rect 255044 396986 255096 396992
rect 254872 396222 254992 396250
rect 254768 393984 254820 393990
rect 254768 393926 254820 393932
rect 254872 393314 254900 396222
rect 254952 396160 255004 396166
rect 254952 396102 255004 396108
rect 254596 393286 254900 393314
rect 254596 351218 254624 393286
rect 254584 351212 254636 351218
rect 254584 351154 254636 351160
rect 254492 24132 254544 24138
rect 254492 24074 254544 24080
rect 254400 17400 254452 17406
rect 254400 17342 254452 17348
rect 254308 17264 254360 17270
rect 254308 17206 254360 17212
rect 254124 6248 254176 6254
rect 254124 6190 254176 6196
rect 254032 6180 254084 6186
rect 254032 6122 254084 6128
rect 254674 5128 254730 5137
rect 254674 5063 254730 5072
rect 251180 4888 251232 4894
rect 251180 4830 251232 4836
rect 252744 4888 252796 4894
rect 252744 4830 252796 4836
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 248420 3528 248472 3534
rect 248420 3470 248472 3476
rect 247604 480 247632 3470
rect 248788 3256 248840 3262
rect 248788 3198 248840 3204
rect 248800 480 248828 3198
rect 249984 3120 250036 3126
rect 249984 3062 250036 3068
rect 249996 480 250024 3062
rect 251192 480 251220 4830
rect 252376 4820 252428 4826
rect 252376 4762 252428 4768
rect 252388 480 252416 4762
rect 253478 3360 253534 3369
rect 253478 3295 253534 3304
rect 253492 480 253520 3295
rect 254688 480 254716 5063
rect 254964 4826 254992 396102
rect 255056 395350 255084 396986
rect 255332 396658 255360 400044
rect 255424 398478 255452 400044
rect 255412 398472 255464 398478
rect 255412 398414 255464 398420
rect 255516 398070 255544 400044
rect 255504 398064 255556 398070
rect 255504 398006 255556 398012
rect 255608 397905 255636 400044
rect 261484 398812 261536 398818
rect 261484 398754 261536 398760
rect 256238 398304 256294 398313
rect 256238 398239 256294 398248
rect 256054 398032 256110 398041
rect 256054 397967 256110 397976
rect 255594 397896 255650 397905
rect 255594 397831 255650 397840
rect 255964 397724 256016 397730
rect 255964 397666 256016 397672
rect 255976 397390 256004 397666
rect 255964 397384 256016 397390
rect 255964 397326 256016 397332
rect 255964 397180 256016 397186
rect 255964 397122 256016 397128
rect 255332 396630 255452 396658
rect 255318 395720 255374 395729
rect 255318 395655 255374 395664
rect 255044 395344 255096 395350
rect 255044 395286 255096 395292
rect 255332 16574 255360 395655
rect 255424 25566 255452 396630
rect 255412 25560 255464 25566
rect 255412 25502 255464 25508
rect 255332 16546 255912 16574
rect 254952 4820 255004 4826
rect 254952 4762 255004 4768
rect 255884 480 255912 16546
rect 255976 3466 256004 397122
rect 256068 6322 256096 397967
rect 256252 397594 256280 398239
rect 256700 398200 256752 398206
rect 256700 398142 256752 398148
rect 256332 397792 256384 397798
rect 256332 397734 256384 397740
rect 256148 397588 256200 397594
rect 256148 397530 256200 397536
rect 256240 397588 256292 397594
rect 256240 397530 256292 397536
rect 256160 397474 256188 397530
rect 256160 397446 256280 397474
rect 256148 397384 256200 397390
rect 256148 397326 256200 397332
rect 256160 14958 256188 397326
rect 256252 60042 256280 397446
rect 256344 60110 256372 397734
rect 256332 60104 256384 60110
rect 256332 60046 256384 60052
rect 256240 60036 256292 60042
rect 256240 59978 256292 59984
rect 256148 14952 256200 14958
rect 256148 14894 256200 14900
rect 256056 6316 256108 6322
rect 256056 6258 256108 6264
rect 255964 3460 256016 3466
rect 255964 3402 256016 3408
rect 228702 354 228814 480
rect 228560 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 398142
rect 258816 398064 258868 398070
rect 258816 398006 258868 398012
rect 257528 397996 257580 398002
rect 257528 397938 257580 397944
rect 257436 397860 257488 397866
rect 257436 397802 257488 397808
rect 257342 396536 257398 396545
rect 257342 396471 257398 396480
rect 257356 3602 257384 396471
rect 257448 8974 257476 397802
rect 257540 304298 257568 397938
rect 258724 397656 258776 397662
rect 258724 397598 258776 397604
rect 258736 333266 258764 397598
rect 258828 334626 258856 398006
rect 258816 334620 258868 334626
rect 258816 334562 258868 334568
rect 258724 333260 258776 333266
rect 258724 333202 258776 333208
rect 257528 304292 257580 304298
rect 257528 304234 257580 304240
rect 261496 180130 261524 398754
rect 264244 398608 264296 398614
rect 264244 398550 264296 398556
rect 262220 354340 262272 354346
rect 262220 354282 262272 354288
rect 261484 180124 261536 180130
rect 261484 180066 261536 180072
rect 262232 16574 262260 354282
rect 264256 28286 264284 398550
rect 264336 398540 264388 398546
rect 264336 398482 264388 398488
rect 264348 182850 264376 398482
rect 264336 182844 264388 182850
rect 264336 182786 264388 182792
rect 265636 86970 265664 444615
rect 265728 299470 265756 444926
rect 265806 443728 265862 443737
rect 265806 443663 265862 443672
rect 265820 404326 265848 443663
rect 265912 431934 265940 445198
rect 265900 431928 265952 431934
rect 265900 431870 265952 431876
rect 267016 426426 267044 445266
rect 273902 444952 273958 444961
rect 273902 444887 273958 444896
rect 269856 444780 269908 444786
rect 269856 444722 269908 444728
rect 268382 444544 268438 444553
rect 268382 444479 268438 444488
rect 267004 426420 267056 426426
rect 267004 426362 267056 426368
rect 265808 404320 265860 404326
rect 265808 404262 265860 404268
rect 266360 395820 266412 395826
rect 266360 395762 266412 395768
rect 265716 299464 265768 299470
rect 265716 299406 265768 299412
rect 265624 86964 265676 86970
rect 265624 86906 265676 86912
rect 264244 28280 264296 28286
rect 264244 28222 264296 28228
rect 266372 16574 266400 395762
rect 268396 126954 268424 444479
rect 269764 398404 269816 398410
rect 269764 398346 269816 398352
rect 269120 395752 269172 395758
rect 269120 395694 269172 395700
rect 268384 126948 268436 126954
rect 268384 126890 268436 126896
rect 269132 16574 269160 395694
rect 269776 29646 269804 398346
rect 269868 206990 269896 444722
rect 271236 444712 271288 444718
rect 271236 444654 271288 444660
rect 271144 398336 271196 398342
rect 271144 398278 271196 398284
rect 269856 206984 269908 206990
rect 269856 206926 269908 206932
rect 271156 31074 271184 398278
rect 271248 193186 271276 444654
rect 273258 354376 273314 354385
rect 273258 354311 273314 354320
rect 271236 193180 271288 193186
rect 271236 193122 271288 193128
rect 271144 31068 271196 31074
rect 271144 31010 271196 31016
rect 269764 29640 269816 29646
rect 269764 29582 269816 29588
rect 271880 17672 271932 17678
rect 271880 17614 271932 17620
rect 271892 16574 271920 17614
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 271892 16546 272472 16574
rect 257436 8968 257488 8974
rect 257436 8910 257488 8916
rect 261760 6044 261812 6050
rect 261760 5986 261812 5992
rect 259460 4140 259512 4146
rect 259460 4082 259512 4088
rect 258264 4072 258316 4078
rect 258264 4014 258316 4020
rect 257344 3596 257396 3602
rect 257344 3538 257396 3544
rect 258276 480 258304 4014
rect 259472 480 259500 4082
rect 260656 4004 260708 4010
rect 260656 3946 260708 3952
rect 260668 480 260696 3946
rect 261772 480 261800 5986
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 265348 6112 265400 6118
rect 265348 6054 265400 6060
rect 264152 3868 264204 3874
rect 264152 3810 264204 3816
rect 264164 480 264192 3810
rect 265360 480 265388 6054
rect 266556 480 266584 16546
rect 267740 6860 267792 6866
rect 267740 6802 267792 6808
rect 267752 480 267780 6802
rect 268844 6792 268896 6798
rect 268844 6734 268896 6740
rect 268856 480 268884 6734
rect 270052 480 270080 16546
rect 271236 3936 271288 3942
rect 271236 3878 271288 3884
rect 271248 480 271276 3878
rect 272444 480 272472 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 354311
rect 273916 60722 273944 444887
rect 273996 444644 274048 444650
rect 273996 444586 274048 444592
rect 274008 167006 274036 444586
rect 275468 443216 275520 443222
rect 275468 443158 275520 443164
rect 275376 443148 275428 443154
rect 275376 443090 275428 443096
rect 275388 398274 275416 443090
rect 274088 398268 274140 398274
rect 274088 398210 274140 398216
rect 275376 398268 275428 398274
rect 275376 398210 275428 398216
rect 274100 184210 274128 398210
rect 275480 398206 275508 443158
rect 293130 442776 293186 442785
rect 293130 442711 293186 442720
rect 292946 442504 293002 442513
rect 292946 442439 293002 442448
rect 292960 401062 292988 442439
rect 292948 401056 293000 401062
rect 292948 400998 293000 401004
rect 293144 400897 293172 442711
rect 293236 400994 293264 449890
rect 293316 448656 293368 448662
rect 293316 448598 293368 448604
rect 293224 400988 293276 400994
rect 293224 400930 293276 400936
rect 293328 400926 293356 448598
rect 293408 448588 293460 448594
rect 293408 448530 293460 448536
rect 293420 401130 293448 448530
rect 296088 447846 296116 458594
rect 297192 449886 297220 525943
rect 297376 524385 297404 600102
rect 297468 598942 297496 631479
rect 297546 628552 297602 628561
rect 297546 628487 297602 628496
rect 297456 598936 297508 598942
rect 297456 598878 297508 598884
rect 297362 524376 297418 524385
rect 297362 524311 297418 524320
rect 297468 521665 297496 598878
rect 297560 598806 297588 628487
rect 297638 608288 297694 608297
rect 297638 608223 297694 608232
rect 297548 598800 297600 598806
rect 297548 598742 297600 598748
rect 297454 521656 297510 521665
rect 297454 521591 297510 521600
rect 297468 509234 297496 521591
rect 297560 518673 297588 598742
rect 297546 518664 297602 518673
rect 297546 518599 297602 518608
rect 297560 517585 297588 518599
rect 297546 517576 297602 517585
rect 297546 517511 297602 517520
rect 297376 509206 297496 509234
rect 297376 488481 297404 509206
rect 297652 498409 297680 608223
rect 297744 523297 297772 633111
rect 297822 630184 297878 630193
rect 297822 630119 297878 630128
rect 297836 538214 297864 630119
rect 297928 600166 297956 634199
rect 297916 600160 297968 600166
rect 297916 600102 297968 600108
rect 298020 598874 298048 636919
rect 298008 598868 298060 598874
rect 298008 598810 298060 598816
rect 298020 598602 298048 598810
rect 298008 598596 298060 598602
rect 298008 598538 298060 598544
rect 317694 597544 317750 597553
rect 317694 597479 317750 597488
rect 320086 597544 320142 597553
rect 320086 597479 320142 597488
rect 320914 597544 320970 597553
rect 320914 597479 320970 597488
rect 322202 597544 322258 597553
rect 322202 597479 322258 597488
rect 322938 597544 322994 597553
rect 322938 597479 322994 597488
rect 324318 597544 324374 597553
rect 324318 597479 324374 597488
rect 326158 597544 326214 597553
rect 326158 597479 326214 597488
rect 329838 597544 329894 597553
rect 329838 597479 329894 597488
rect 345018 597544 345074 597553
rect 345018 597479 345074 597488
rect 360198 597544 360254 597553
rect 360198 597479 360254 597488
rect 313278 597272 313334 597281
rect 313278 597207 313334 597216
rect 313292 596902 313320 597207
rect 299296 596896 299348 596902
rect 299296 596838 299348 596844
rect 313280 596896 313332 596902
rect 313280 596838 313332 596844
rect 314658 596864 314714 596873
rect 299204 596828 299256 596834
rect 299204 596770 299256 596776
rect 298744 584452 298796 584458
rect 298744 584394 298796 584400
rect 297836 538186 297956 538214
rect 297822 524376 297878 524385
rect 297822 524311 297878 524320
rect 297730 523288 297786 523297
rect 297730 523223 297786 523232
rect 297638 498400 297694 498409
rect 297638 498335 297694 498344
rect 297456 489864 297508 489870
rect 297456 489806 297508 489812
rect 297362 488472 297418 488481
rect 297362 488407 297418 488416
rect 297362 488336 297418 488345
rect 297362 488271 297418 488280
rect 297180 449880 297232 449886
rect 297180 449822 297232 449828
rect 297376 448458 297404 488271
rect 297364 448452 297416 448458
rect 297364 448394 297416 448400
rect 297468 448322 297496 489806
rect 297548 488504 297600 488510
rect 297548 488446 297600 488452
rect 297560 488170 297588 488446
rect 297652 488442 297680 498335
rect 297744 489870 297772 523223
rect 297836 518894 297864 524311
rect 297928 521914 297956 538186
rect 298006 527096 298062 527105
rect 298006 527031 298062 527040
rect 298020 526794 298048 527031
rect 298008 526788 298060 526794
rect 298008 526730 298060 526736
rect 297928 521886 298048 521914
rect 298020 520305 298048 521886
rect 298006 520296 298062 520305
rect 298006 520231 298062 520240
rect 297836 518866 297956 518894
rect 297824 498840 297876 498846
rect 297824 498782 297876 498788
rect 297836 498681 297864 498782
rect 297822 498672 297878 498681
rect 297822 498607 297878 498616
rect 297732 489864 297784 489870
rect 297928 489841 297956 518866
rect 297732 489806 297784 489812
rect 297914 489832 297970 489841
rect 297914 489767 297970 489776
rect 297732 488504 297784 488510
rect 297732 488446 297784 488452
rect 297822 488472 297878 488481
rect 297640 488436 297692 488442
rect 297640 488378 297692 488384
rect 297548 488164 297600 488170
rect 297548 488106 297600 488112
rect 297456 448316 297508 448322
rect 297456 448258 297508 448264
rect 297560 448254 297588 488106
rect 297638 452432 297694 452441
rect 297638 452367 297694 452376
rect 297652 451314 297680 452367
rect 297640 451308 297692 451314
rect 297640 451250 297692 451256
rect 297744 448526 297772 488446
rect 297822 488407 297878 488416
rect 297732 448520 297784 448526
rect 297732 448462 297784 448468
rect 297836 448390 297864 488407
rect 297928 449857 297956 489767
rect 298020 488510 298048 520231
rect 298008 488504 298060 488510
rect 298008 488446 298060 488452
rect 298020 488374 298048 488446
rect 298008 488368 298060 488374
rect 298008 488310 298060 488316
rect 298100 488300 298152 488306
rect 298100 488242 298152 488248
rect 298112 487830 298140 488242
rect 298100 487824 298152 487830
rect 298100 487766 298152 487772
rect 298008 458448 298060 458454
rect 298008 458390 298060 458396
rect 298020 450770 298048 458390
rect 298008 450764 298060 450770
rect 298008 450706 298060 450712
rect 297914 449848 297970 449857
rect 297914 449783 297970 449792
rect 297824 448384 297876 448390
rect 297824 448326 297876 448332
rect 298006 448352 298062 448361
rect 298006 448287 298062 448296
rect 297548 448248 297600 448254
rect 297548 448190 297600 448196
rect 296076 447840 296128 447846
rect 296076 447782 296128 447788
rect 298020 447574 298048 448287
rect 298008 447568 298060 447574
rect 298008 447510 298060 447516
rect 296352 447500 296404 447506
rect 296352 447442 296404 447448
rect 296168 447296 296220 447302
rect 295982 447264 296038 447273
rect 296168 447238 296220 447244
rect 295982 447199 296038 447208
rect 293868 445188 293920 445194
rect 293868 445130 293920 445136
rect 293684 445120 293736 445126
rect 293684 445062 293736 445068
rect 293592 444916 293644 444922
rect 293592 444858 293644 444864
rect 293500 444848 293552 444854
rect 293500 444790 293552 444796
rect 293408 401124 293460 401130
rect 293408 401066 293460 401072
rect 293316 400920 293368 400926
rect 293130 400888 293186 400897
rect 293316 400862 293368 400868
rect 293130 400823 293186 400832
rect 293512 398478 293540 444790
rect 293604 398818 293632 444858
rect 293592 398812 293644 398818
rect 293592 398754 293644 398760
rect 293696 398682 293724 445062
rect 293774 442640 293830 442649
rect 293774 442575 293830 442584
rect 293684 398676 293736 398682
rect 293684 398618 293736 398624
rect 293788 398614 293816 442575
rect 293880 401606 293908 445130
rect 295892 444508 295944 444514
rect 295892 444450 295944 444456
rect 295800 444032 295852 444038
rect 295800 443974 295852 443980
rect 293868 401600 293920 401606
rect 293868 401542 293920 401548
rect 293776 398608 293828 398614
rect 293776 398550 293828 398556
rect 295812 398546 295840 443974
rect 295800 398540 295852 398546
rect 295800 398482 295852 398488
rect 278044 398472 278096 398478
rect 278044 398414 278096 398420
rect 293500 398472 293552 398478
rect 293500 398414 293552 398420
rect 275468 398200 275520 398206
rect 275468 398142 275520 398148
rect 275282 397896 275338 397905
rect 275282 397831 275338 397840
rect 275296 185638 275324 397831
rect 276020 395684 276072 395690
rect 276020 395626 276072 395632
rect 275284 185632 275336 185638
rect 275284 185574 275336 185580
rect 274088 184204 274140 184210
rect 274088 184146 274140 184152
rect 273996 167000 274048 167006
rect 273996 166942 274048 166948
rect 273904 60716 273956 60722
rect 273904 60658 273956 60664
rect 276032 16574 276060 395626
rect 277400 392828 277452 392834
rect 277400 392770 277452 392776
rect 277412 16574 277440 392770
rect 278056 82142 278084 398414
rect 293960 395616 294012 395622
rect 291198 395584 291254 395593
rect 293960 395558 294012 395564
rect 291198 395519 291254 395528
rect 281540 392760 281592 392766
rect 281540 392702 281592 392708
rect 278044 82136 278096 82142
rect 278044 82078 278096 82084
rect 280160 25968 280212 25974
rect 280160 25910 280212 25916
rect 278780 17604 278832 17610
rect 278780 17546 278832 17552
rect 278792 16574 278820 17546
rect 280172 16574 280200 25910
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276018 6760 276074 6769
rect 276018 6695 276074 6704
rect 274822 3224 274878 3233
rect 274822 3159 274878 3168
rect 274836 480 274864 3159
rect 276032 480 276060 6695
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 392702
rect 284300 355496 284352 355502
rect 284300 355438 284352 355444
rect 282920 17536 282972 17542
rect 282920 17478 282972 17484
rect 282932 16574 282960 17478
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 3874 284340 355438
rect 288440 87848 288492 87854
rect 288440 87790 288492 87796
rect 284392 25900 284444 25906
rect 284392 25842 284444 25848
rect 284300 3868 284352 3874
rect 284300 3810 284352 3816
rect 284404 3482 284432 25842
rect 287060 25832 287112 25838
rect 287060 25774 287112 25780
rect 285680 18964 285732 18970
rect 285680 18906 285732 18912
rect 285692 16574 285720 18906
rect 287072 16574 287100 25774
rect 288452 16574 288480 87790
rect 289818 18864 289874 18873
rect 289818 18799 289874 18808
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 285036 3868 285088 3874
rect 285036 3810 285088 3816
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3810
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 18799
rect 291212 16574 291240 395519
rect 292578 18728 292634 18737
rect 292578 18663 292634 18672
rect 292592 16574 292620 18663
rect 293972 16574 294000 395558
rect 295904 365702 295932 444450
rect 295892 365696 295944 365702
rect 295892 365638 295944 365644
rect 295996 139398 296024 447199
rect 296074 442368 296130 442377
rect 296074 442303 296130 442312
rect 295984 139392 296036 139398
rect 295984 139334 296036 139340
rect 296088 100706 296116 442303
rect 296180 179382 296208 447238
rect 296260 447228 296312 447234
rect 296260 447170 296312 447176
rect 296272 219434 296300 447170
rect 296364 259418 296392 447442
rect 296628 447432 296680 447438
rect 296628 447374 296680 447380
rect 296444 447364 296496 447370
rect 296444 447306 296496 447312
rect 296456 273222 296484 447306
rect 296536 446276 296588 446282
rect 296536 446218 296588 446224
rect 296548 313274 296576 446218
rect 296640 325650 296668 447374
rect 298756 446418 298784 584394
rect 299216 488238 299244 596770
rect 299308 488306 299336 596838
rect 314658 596799 314660 596808
rect 314712 596799 314714 596808
rect 314660 596770 314712 596776
rect 317708 596766 317736 597479
rect 319994 597408 320050 597417
rect 319994 597343 320050 597352
rect 320008 597310 320036 597343
rect 319996 597304 320048 597310
rect 319996 597246 320048 597252
rect 318708 597168 318760 597174
rect 318708 597110 318760 597116
rect 318720 596766 318748 597110
rect 317696 596760 317748 596766
rect 317696 596702 317748 596708
rect 318708 596760 318760 596766
rect 318708 596702 318760 596708
rect 311898 596592 311954 596601
rect 311898 596527 311954 596536
rect 311912 596222 311940 596527
rect 320008 596494 320036 597246
rect 320100 596698 320128 597479
rect 320928 596970 320956 597479
rect 320916 596964 320968 596970
rect 320916 596906 320968 596912
rect 320088 596692 320140 596698
rect 320088 596634 320140 596640
rect 320928 596630 320956 596906
rect 320916 596624 320968 596630
rect 320916 596566 320968 596572
rect 322216 596562 322244 597479
rect 322952 597038 322980 597479
rect 322940 597032 322992 597038
rect 322940 596974 322992 596980
rect 322204 596556 322256 596562
rect 322204 596498 322256 596504
rect 319996 596488 320048 596494
rect 319996 596430 320048 596436
rect 322952 596426 322980 596974
rect 322940 596420 322992 596426
rect 322940 596362 322992 596368
rect 299388 596216 299440 596222
rect 299388 596158 299440 596164
rect 311900 596216 311952 596222
rect 311900 596158 311952 596164
rect 299296 488300 299348 488306
rect 299296 488242 299348 488248
rect 299204 488232 299256 488238
rect 299204 488174 299256 488180
rect 299400 487150 299428 596158
rect 324332 587246 324360 597479
rect 324410 597408 324466 597417
rect 324410 597343 324466 597352
rect 324424 597106 324452 597343
rect 326172 597242 326200 597479
rect 326160 597236 326212 597242
rect 326160 597178 326212 597184
rect 324412 597100 324464 597106
rect 324412 597042 324464 597048
rect 324424 596358 324452 597042
rect 324412 596352 324464 596358
rect 324412 596294 324464 596300
rect 326172 596290 326200 597178
rect 326160 596284 326212 596290
rect 326160 596226 326212 596232
rect 329852 589966 329880 597479
rect 335358 597408 335414 597417
rect 335358 597343 335360 597352
rect 335412 597343 335414 597352
rect 335360 597314 335412 597320
rect 339498 597000 339554 597009
rect 339498 596935 339554 596944
rect 329840 589960 329892 589966
rect 329840 589902 329892 589908
rect 339512 588606 339540 596935
rect 339500 588600 339552 588606
rect 339500 588542 339552 588548
rect 324320 587240 324372 587246
rect 324320 587182 324372 587188
rect 345032 581670 345060 597479
rect 349158 597136 349214 597145
rect 349158 597071 349214 597080
rect 349172 583030 349200 597071
rect 354678 596320 354734 596329
rect 354678 596255 354734 596264
rect 354692 584458 354720 596255
rect 360212 585886 360240 597479
rect 360200 585880 360252 585886
rect 360200 585822 360252 585828
rect 354680 584452 354732 584458
rect 354680 584394 354732 584400
rect 349160 583024 349212 583030
rect 349160 582966 349212 582972
rect 345020 581664 345072 581670
rect 345020 581606 345072 581612
rect 314290 488472 314346 488481
rect 314290 488407 314346 488416
rect 315394 488472 315450 488481
rect 315394 488407 315450 488416
rect 314304 488306 314332 488407
rect 314292 488300 314344 488306
rect 314292 488242 314344 488248
rect 315408 488238 315436 488407
rect 315396 488232 315448 488238
rect 315396 488174 315448 488180
rect 313002 487928 313058 487937
rect 313002 487863 313058 487872
rect 324410 487928 324466 487937
rect 324410 487863 324466 487872
rect 313016 487830 313044 487863
rect 312544 487824 312596 487830
rect 312544 487766 312596 487772
rect 313004 487824 313056 487830
rect 313004 487766 313056 487772
rect 312556 487150 312584 487766
rect 319444 487620 319496 487626
rect 319444 487562 319496 487568
rect 318064 487552 318116 487558
rect 318064 487494 318116 487500
rect 318076 487257 318104 487494
rect 319456 487257 319484 487562
rect 319994 487520 320050 487529
rect 319994 487455 319996 487464
rect 320048 487455 320050 487464
rect 322938 487520 322994 487529
rect 322938 487455 322994 487464
rect 319996 487426 320048 487432
rect 318062 487248 318118 487257
rect 318062 487183 318118 487192
rect 319442 487248 319498 487257
rect 319442 487183 319498 487192
rect 299388 487144 299440 487150
rect 299388 487086 299440 487092
rect 311900 487144 311952 487150
rect 311900 487086 311952 487092
rect 312544 487144 312596 487150
rect 312544 487086 312596 487092
rect 311912 464506 311940 487086
rect 318076 475522 318104 487183
rect 318064 475516 318116 475522
rect 318064 475458 318116 475464
rect 319456 473346 319484 487183
rect 320008 485246 320036 487426
rect 322952 487422 322980 487455
rect 322940 487416 322992 487422
rect 322202 487384 322258 487393
rect 322940 487358 322992 487364
rect 322202 487319 322258 487328
rect 322216 487286 322244 487319
rect 322204 487280 322256 487286
rect 320822 487248 320878 487257
rect 322204 487222 322256 487228
rect 320822 487183 320824 487192
rect 320876 487183 320878 487192
rect 320824 487154 320876 487160
rect 319996 485240 320048 485246
rect 319996 485182 320048 485188
rect 320836 479602 320864 487154
rect 320824 479596 320876 479602
rect 320824 479538 320876 479544
rect 322216 474706 322244 487222
rect 322952 481098 322980 487358
rect 324424 487354 324452 487863
rect 326618 487792 326674 487801
rect 326618 487727 326674 487736
rect 326632 487694 326660 487727
rect 326620 487688 326672 487694
rect 326620 487630 326672 487636
rect 324412 487348 324464 487354
rect 324412 487290 324464 487296
rect 324318 487248 324374 487257
rect 324318 487183 324374 487192
rect 322940 481092 322992 481098
rect 322940 481034 322992 481040
rect 322204 474700 322256 474706
rect 322204 474642 322256 474648
rect 319444 473340 319496 473346
rect 319444 473282 319496 473288
rect 324332 472734 324360 487183
rect 324424 486606 324452 487290
rect 324412 486600 324464 486606
rect 324412 486542 324464 486548
rect 326632 484362 326660 487630
rect 329838 487248 329894 487257
rect 329838 487183 329894 487192
rect 335358 487248 335414 487257
rect 335358 487183 335414 487192
rect 339498 487248 339554 487257
rect 339498 487183 339554 487192
rect 345018 487248 345074 487257
rect 345018 487183 345074 487192
rect 349158 487248 349214 487257
rect 349158 487183 349214 487192
rect 354678 487248 354734 487257
rect 354678 487183 354734 487192
rect 360198 487248 360254 487257
rect 360198 487183 360254 487192
rect 326620 484356 326672 484362
rect 326620 484298 326672 484304
rect 329852 475454 329880 487183
rect 329840 475448 329892 475454
rect 329840 475390 329892 475396
rect 335372 474094 335400 487183
rect 339512 479670 339540 487183
rect 339500 479664 339552 479670
rect 339500 479606 339552 479612
rect 335360 474088 335412 474094
rect 335360 474030 335412 474036
rect 324320 472728 324372 472734
rect 324320 472670 324372 472676
rect 311900 464500 311952 464506
rect 311900 464442 311952 464448
rect 345032 463146 345060 487183
rect 345020 463140 345072 463146
rect 345020 463082 345072 463088
rect 349172 461718 349200 487183
rect 354692 478242 354720 487183
rect 360212 481030 360240 487183
rect 360200 481024 360252 481030
rect 360200 480966 360252 480972
rect 354680 478236 354732 478242
rect 354680 478178 354732 478184
rect 395356 478174 395384 699654
rect 395344 478168 395396 478174
rect 395344 478110 395396 478116
rect 399496 468586 399524 700334
rect 403636 476882 403664 700402
rect 405016 489190 405044 700538
rect 429856 700534 429884 703520
rect 409144 700528 409196 700534
rect 409144 700470 409196 700476
rect 429844 700528 429896 700534
rect 429844 700470 429896 700476
rect 406384 700324 406436 700330
rect 406384 700266 406436 700272
rect 405004 489184 405056 489190
rect 405004 489126 405056 489132
rect 403624 476876 403676 476882
rect 403624 476818 403676 476824
rect 399484 468580 399536 468586
rect 399484 468522 399536 468528
rect 406396 465798 406424 700266
rect 407946 636440 408002 636449
rect 407946 636375 408002 636384
rect 407670 635352 407726 635361
rect 407670 635287 407726 635296
rect 407578 628008 407634 628017
rect 407578 627943 407634 627952
rect 407592 598806 407620 627943
rect 407580 598800 407632 598806
rect 407580 598742 407632 598748
rect 406476 596352 406528 596358
rect 406476 596294 406528 596300
rect 406384 465792 406436 465798
rect 406384 465734 406436 465740
rect 349160 461712 349212 461718
rect 349160 461654 349212 461660
rect 406488 460290 406516 596294
rect 407684 585818 407712 635287
rect 407762 629640 407818 629649
rect 407762 629575 407818 629584
rect 407672 585812 407724 585818
rect 407672 585754 407724 585760
rect 407684 526561 407712 585754
rect 407670 526552 407726 526561
rect 407670 526487 407726 526496
rect 407670 523288 407726 523297
rect 407670 523223 407726 523232
rect 407578 520976 407634 520985
rect 407578 520911 407634 520920
rect 407394 517984 407450 517993
rect 407394 517919 407450 517928
rect 407408 488209 407436 517919
rect 407592 488345 407620 520911
rect 407684 489870 407712 523223
rect 407776 520305 407804 629575
rect 407854 607744 407910 607753
rect 407854 607679 407910 607688
rect 407762 520296 407818 520305
rect 407762 520231 407818 520240
rect 407672 489864 407724 489870
rect 407672 489806 407724 489812
rect 407776 488374 407804 520231
rect 407868 498409 407896 607679
rect 407960 598874 407988 636375
rect 408130 633720 408186 633729
rect 408130 633655 408186 633664
rect 408038 632632 408094 632641
rect 408038 632567 408094 632576
rect 407948 598868 408000 598874
rect 407948 598810 408000 598816
rect 407948 596556 408000 596562
rect 407948 596498 408000 596504
rect 407854 498400 407910 498409
rect 407854 498335 407910 498344
rect 407868 488442 407896 498335
rect 407856 488436 407908 488442
rect 407856 488378 407908 488384
rect 407960 488374 407988 596498
rect 408052 523297 408080 632567
rect 408144 600030 408172 633655
rect 408222 631000 408278 631009
rect 408222 630935 408278 630944
rect 408132 600024 408184 600030
rect 408132 599966 408184 599972
rect 408236 598942 408264 630935
rect 408314 610056 408370 610065
rect 408314 609991 408370 610000
rect 408224 598936 408276 598942
rect 408224 598878 408276 598884
rect 408132 596488 408184 596494
rect 408132 596430 408184 596436
rect 408038 523288 408094 523297
rect 408038 523223 408094 523232
rect 408038 498264 408094 498273
rect 408038 498199 408094 498208
rect 407764 488368 407816 488374
rect 407578 488336 407634 488345
rect 407764 488310 407816 488316
rect 407948 488368 408000 488374
rect 407948 488310 408000 488316
rect 407578 488271 407634 488280
rect 407394 488200 407450 488209
rect 407394 488135 407450 488144
rect 407960 487830 407988 488310
rect 407948 487824 408000 487830
rect 407948 487766 408000 487772
rect 408052 463078 408080 498199
rect 408144 488442 408172 596430
rect 408224 596420 408276 596426
rect 408224 596362 408276 596368
rect 408236 488510 408264 596362
rect 408328 500313 408356 609991
rect 408406 608696 408462 608705
rect 408406 608631 408462 608640
rect 408314 500304 408370 500313
rect 408314 500239 408370 500248
rect 408224 488504 408276 488510
rect 408224 488446 408276 488452
rect 408132 488436 408184 488442
rect 408132 488378 408184 488384
rect 408144 488306 408172 488378
rect 408132 488300 408184 488306
rect 408132 488242 408184 488248
rect 408236 488238 408264 488446
rect 408224 488232 408276 488238
rect 408224 488174 408276 488180
rect 408328 488170 408356 500239
rect 408420 498681 408448 608631
rect 408406 498672 408462 498681
rect 408406 498607 408462 498616
rect 408420 498273 408448 498607
rect 408406 498264 408462 498273
rect 408406 498199 408462 498208
rect 408316 488164 408368 488170
rect 408316 488106 408368 488112
rect 409156 467226 409184 700470
rect 462332 700466 462360 703520
rect 462320 700460 462372 700466
rect 462320 700402 462372 700408
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 509884 700324 509936 700330
rect 509884 700266 509936 700272
rect 508504 670744 508556 670750
rect 508504 670686 508556 670692
rect 501604 630692 501656 630698
rect 501604 630634 501656 630640
rect 440238 597544 440294 597553
rect 440238 597479 440294 597488
rect 449898 597544 449954 597553
rect 449898 597479 449954 597488
rect 459558 597544 459614 597553
rect 459558 597479 459614 597488
rect 427818 597408 427874 597417
rect 427818 597343 427874 597352
rect 430578 597408 430634 597417
rect 430578 597343 430634 597352
rect 434718 597408 434774 597417
rect 434718 597343 434774 597352
rect 427832 597310 427860 597343
rect 427820 597304 427872 597310
rect 422574 597272 422630 597281
rect 422574 597207 422630 597216
rect 426438 597272 426494 597281
rect 427820 597246 427872 597252
rect 426438 597207 426494 597216
rect 409326 596864 409382 596873
rect 409326 596799 409382 596808
rect 409236 596216 409288 596222
rect 409236 596158 409288 596164
rect 409248 483750 409276 596158
rect 409340 485110 409368 596799
rect 422588 596562 422616 597207
rect 426452 597174 426480 597207
rect 426440 597168 426492 597174
rect 426440 597110 426492 597116
rect 423678 597000 423734 597009
rect 423678 596935 423734 596944
rect 429198 597000 429254 597009
rect 430592 596970 430620 597343
rect 434732 597242 434760 597343
rect 434720 597236 434772 597242
rect 434720 597178 434772 597184
rect 433338 597136 433394 597145
rect 433338 597071 433394 597080
rect 434718 597136 434774 597145
rect 434718 597071 434720 597080
rect 433352 597038 433380 597071
rect 434772 597071 434774 597080
rect 434720 597042 434772 597048
rect 433340 597032 433392 597038
rect 431958 597000 432014 597009
rect 429198 596935 429254 596944
rect 430580 596964 430632 596970
rect 422576 596556 422628 596562
rect 422576 596498 422628 596504
rect 423692 596494 423720 596935
rect 429212 596902 429240 596935
rect 433340 596974 433392 596980
rect 431958 596935 432014 596944
rect 430580 596906 430632 596912
rect 429200 596896 429252 596902
rect 429200 596838 429252 596844
rect 431972 596834 432000 596935
rect 431960 596828 432012 596834
rect 431960 596770 432012 596776
rect 434718 596728 434774 596737
rect 434718 596663 434774 596672
rect 423680 596488 423732 596494
rect 423680 596430 423732 596436
rect 425058 596456 425114 596465
rect 425058 596391 425060 596400
rect 425112 596391 425114 596400
rect 425060 596362 425112 596368
rect 434732 596358 434760 596663
rect 434720 596352 434772 596358
rect 434720 596294 434772 596300
rect 409420 596284 409472 596290
rect 409420 596226 409472 596232
rect 409432 486538 409460 596226
rect 440252 592686 440280 597479
rect 444378 596728 444434 596737
rect 444378 596663 444434 596672
rect 444392 596290 444420 596663
rect 444380 596284 444432 596290
rect 444380 596226 444432 596232
rect 440240 592680 440292 592686
rect 440240 592622 440292 592628
rect 449912 587178 449940 597479
rect 455418 596320 455474 596329
rect 455418 596255 455474 596264
rect 455432 596222 455460 596255
rect 455420 596216 455472 596222
rect 455420 596158 455472 596164
rect 449900 587172 449952 587178
rect 449900 587114 449952 587120
rect 459572 580310 459600 597479
rect 470598 596320 470654 596329
rect 470598 596255 470654 596264
rect 470612 589937 470640 596255
rect 470598 589928 470654 589937
rect 470598 589863 470654 589872
rect 459560 580304 459612 580310
rect 459560 580246 459612 580252
rect 425060 488504 425112 488510
rect 422574 488472 422630 488481
rect 422574 488407 422630 488416
rect 423678 488472 423734 488481
rect 423678 488407 423680 488416
rect 422588 488374 422616 488407
rect 423732 488407 423734 488416
rect 425058 488472 425060 488481
rect 425112 488472 425114 488481
rect 425058 488407 425114 488416
rect 423680 488378 423732 488384
rect 422576 488368 422628 488374
rect 422576 488310 422628 488316
rect 465078 488336 465134 488345
rect 465078 488271 465134 488280
rect 429198 488200 429254 488209
rect 429198 488135 429254 488144
rect 434718 488200 434774 488209
rect 434718 488135 434774 488144
rect 426438 487656 426494 487665
rect 426438 487591 426494 487600
rect 427818 487656 427874 487665
rect 427818 487591 427820 487600
rect 426452 487558 426480 487591
rect 427872 487591 427874 487600
rect 427820 487562 427872 487568
rect 426440 487552 426492 487558
rect 426440 487494 426492 487500
rect 429212 487490 429240 488135
rect 430578 487792 430634 487801
rect 430578 487727 430634 487736
rect 429200 487484 429252 487490
rect 429200 487426 429252 487432
rect 430592 487218 430620 487727
rect 434732 487694 434760 488135
rect 434720 487688 434772 487694
rect 434720 487630 434772 487636
rect 433338 487520 433394 487529
rect 433338 487455 433394 487464
rect 433352 487422 433380 487455
rect 433340 487416 433392 487422
rect 432142 487384 432198 487393
rect 433340 487358 433392 487364
rect 434718 487384 434774 487393
rect 432142 487319 432198 487328
rect 434718 487319 434720 487328
rect 432156 487286 432184 487319
rect 434772 487319 434774 487328
rect 434720 487290 434772 487296
rect 432144 487280 432196 487286
rect 432144 487222 432196 487228
rect 434718 487248 434774 487257
rect 430580 487212 430632 487218
rect 440238 487248 440294 487257
rect 434718 487183 434774 487192
rect 436744 487212 436796 487218
rect 430580 487154 430632 487160
rect 409420 486532 409472 486538
rect 409420 486474 409472 486480
rect 409328 485104 409380 485110
rect 409328 485046 409380 485052
rect 409236 483744 409288 483750
rect 409236 483686 409288 483692
rect 434732 482390 434760 487183
rect 440238 487183 440294 487192
rect 444378 487248 444434 487257
rect 444378 487183 444434 487192
rect 449898 487248 449954 487257
rect 449898 487183 449954 487192
rect 455418 487248 455474 487257
rect 455418 487183 455474 487192
rect 459558 487248 459614 487257
rect 465092 487218 465120 488271
rect 470598 487248 470654 487257
rect 459558 487183 459614 487192
rect 465080 487212 465132 487218
rect 436744 487154 436796 487160
rect 434720 482384 434772 482390
rect 434720 482326 434772 482332
rect 409144 467220 409196 467226
rect 409144 467162 409196 467168
rect 436756 465730 436784 487154
rect 440252 471306 440280 487183
rect 440240 471300 440292 471306
rect 440240 471242 440292 471248
rect 436744 465724 436796 465730
rect 436744 465666 436796 465672
rect 444392 464438 444420 487183
rect 449912 468518 449940 487183
rect 455432 469946 455460 487183
rect 459572 476814 459600 487183
rect 470598 487183 470654 487192
rect 465080 487154 465132 487160
rect 459560 476808 459612 476814
rect 459560 476750 459612 476756
rect 455420 469940 455472 469946
rect 455420 469882 455472 469888
rect 449900 468512 449952 468518
rect 449900 468454 449952 468460
rect 470612 467158 470640 487183
rect 501616 482322 501644 630634
rect 504364 616888 504416 616894
rect 504364 616830 504416 616836
rect 502984 510672 503036 510678
rect 502984 510614 503036 510620
rect 501604 482316 501656 482322
rect 501604 482258 501656 482264
rect 470600 467152 470652 467158
rect 470600 467094 470652 467100
rect 444380 464432 444432 464438
rect 444380 464374 444432 464380
rect 408040 463072 408092 463078
rect 408040 463014 408092 463020
rect 406476 460284 406528 460290
rect 406476 460226 406528 460232
rect 502996 460222 503024 510614
rect 504376 464370 504404 616830
rect 507124 563100 507176 563106
rect 507124 563042 507176 563048
rect 504364 464364 504416 464370
rect 504364 464306 504416 464312
rect 507136 461650 507164 563042
rect 508516 463010 508544 670686
rect 509896 469878 509924 700266
rect 512644 643136 512696 643142
rect 512644 643078 512696 643084
rect 511264 536852 511316 536858
rect 511264 536794 511316 536800
rect 511276 472666 511304 536794
rect 512656 474026 512684 643078
rect 516784 576904 516836 576910
rect 516784 576846 516836 576852
rect 514024 524476 514076 524482
rect 514024 524418 514076 524424
rect 514036 479534 514064 524418
rect 516796 480962 516824 576846
rect 516784 480956 516836 480962
rect 516784 480898 516836 480904
rect 514024 479528 514076 479534
rect 514024 479470 514076 479476
rect 527192 475386 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 486470 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 542360 486464 542412 486470
rect 542360 486406 542412 486412
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 483682 580304 683839
rect 580264 483676 580316 483682
rect 580264 483618 580316 483624
rect 527180 475380 527232 475386
rect 527180 475322 527232 475328
rect 512644 474020 512696 474026
rect 512644 473962 512696 473968
rect 511264 472660 511316 472666
rect 511264 472602 511316 472608
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 509884 469872 509936 469878
rect 509884 469814 509936 469820
rect 508504 463004 508556 463010
rect 508504 462946 508556 462952
rect 507124 461644 507176 461650
rect 507124 461586 507176 461592
rect 502984 460216 503036 460222
rect 502984 460158 503036 460164
rect 299664 458992 299716 458998
rect 299664 458934 299716 458940
rect 321284 458992 321336 458998
rect 321284 458934 321336 458940
rect 299388 458788 299440 458794
rect 299388 458730 299440 458736
rect 298928 458516 298980 458522
rect 298928 458458 298980 458464
rect 298836 455660 298888 455666
rect 298836 455602 298888 455608
rect 298848 449206 298876 455602
rect 298940 449274 298968 458458
rect 299020 456816 299072 456822
rect 299020 456758 299072 456764
rect 299032 453354 299060 456758
rect 299020 453348 299072 453354
rect 299020 453290 299072 453296
rect 299400 451994 299428 458730
rect 299480 458720 299532 458726
rect 299480 458662 299532 458668
rect 299492 454782 299520 458662
rect 299572 458584 299624 458590
rect 299572 458526 299624 458532
rect 299584 454850 299612 458526
rect 299572 454844 299624 454850
rect 299572 454786 299624 454792
rect 299480 454776 299532 454782
rect 299480 454718 299532 454724
rect 299388 451988 299440 451994
rect 299388 451930 299440 451936
rect 299676 451274 299704 458934
rect 309048 458312 309100 458318
rect 309048 458254 309100 458260
rect 299756 456068 299808 456074
rect 299756 456010 299808 456016
rect 300768 456068 300820 456074
rect 300768 456010 300820 456016
rect 299768 453506 299796 456010
rect 300320 455666 300702 455682
rect 300780 455666 300808 456010
rect 309060 455940 309088 458254
rect 317420 457292 317472 457298
rect 317420 457234 317472 457240
rect 312636 456000 312688 456006
rect 312688 455948 312938 455954
rect 312636 455942 312938 455948
rect 312648 455926 312938 455942
rect 317432 455940 317460 457234
rect 321296 455940 321324 458934
rect 371516 458924 371568 458930
rect 371516 458866 371568 458872
rect 329656 458788 329708 458794
rect 329656 458730 329708 458736
rect 325792 457224 325844 457230
rect 325792 457166 325844 457172
rect 325804 455940 325832 457166
rect 329668 455940 329696 458730
rect 342536 458720 342588 458726
rect 342536 458662 342588 458668
rect 338028 457156 338080 457162
rect 338028 457098 338080 457104
rect 334164 457088 334216 457094
rect 334164 457030 334216 457036
rect 334176 455940 334204 457030
rect 338040 455940 338068 457098
rect 342548 455940 342576 458662
rect 346400 458652 346452 458658
rect 346400 458594 346452 458600
rect 346412 455940 346440 458594
rect 350908 458584 350960 458590
rect 350908 458526 350960 458532
rect 350920 455940 350948 458526
rect 359280 458516 359332 458522
rect 359280 458458 359332 458464
rect 355968 458244 356020 458250
rect 355968 458186 356020 458192
rect 355980 457502 356008 458186
rect 355968 457496 356020 457502
rect 355968 457438 356020 457444
rect 354772 457020 354824 457026
rect 354772 456962 354824 456968
rect 354784 455940 354812 456962
rect 359292 455940 359320 458458
rect 367652 458448 367704 458454
rect 367652 458390 367704 458396
rect 363144 458380 363196 458386
rect 363144 458322 363196 458328
rect 363156 455940 363184 458322
rect 367664 455940 367692 458390
rect 371528 455940 371556 458866
rect 379888 458856 379940 458862
rect 379888 458798 379940 458804
rect 376024 458244 376076 458250
rect 376024 458186 376076 458192
rect 376036 455940 376064 458186
rect 379900 455940 379928 458798
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 383752 456952 383804 456958
rect 383752 456894 383804 456900
rect 383764 455940 383792 456894
rect 385316 456884 385368 456890
rect 385316 456826 385368 456832
rect 385132 455932 385184 455938
rect 385132 455874 385184 455880
rect 384120 455796 384172 455802
rect 384120 455738 384172 455744
rect 300308 455660 300702 455666
rect 300360 455654 300702 455660
rect 300768 455660 300820 455666
rect 300308 455602 300360 455608
rect 300768 455602 300820 455608
rect 384028 455592 384080 455598
rect 304184 455518 304566 455546
rect 384028 455534 384080 455540
rect 304184 455394 304212 455518
rect 299848 455388 299900 455394
rect 299848 455330 299900 455336
rect 304172 455388 304224 455394
rect 304172 455330 304224 455336
rect 299860 454918 299888 455330
rect 299848 454912 299900 454918
rect 299848 454854 299900 454860
rect 383934 454064 383990 454073
rect 383856 454022 383934 454050
rect 299768 453478 299888 453506
rect 299676 451246 299796 451274
rect 299768 450702 299796 451246
rect 299756 450696 299808 450702
rect 299756 450638 299808 450644
rect 298928 449268 298980 449274
rect 298928 449210 298980 449216
rect 298836 449200 298888 449206
rect 298836 449142 298888 449148
rect 299386 448624 299442 448633
rect 299386 448559 299442 448568
rect 299204 447160 299256 447166
rect 299204 447102 299256 447108
rect 298744 446412 298796 446418
rect 298744 446354 298796 446360
rect 299020 446344 299072 446350
rect 298834 446312 298890 446321
rect 299020 446286 299072 446292
rect 298834 446247 298890 446256
rect 298560 446208 298612 446214
rect 298560 446150 298612 446156
rect 297456 443964 297508 443970
rect 297456 443906 297508 443912
rect 296904 443828 296956 443834
rect 296904 443770 296956 443776
rect 296812 443080 296864 443086
rect 296812 443022 296864 443028
rect 296824 439521 296852 443022
rect 296810 439512 296866 439521
rect 296810 439447 296866 439456
rect 296916 434761 296944 443770
rect 297364 443760 297416 443766
rect 297364 443702 297416 443708
rect 296902 434752 296958 434761
rect 296902 434687 296958 434696
rect 297376 408241 297404 443702
rect 297468 413001 297496 443906
rect 297640 443896 297692 443902
rect 297640 443838 297692 443844
rect 297548 443692 297600 443698
rect 297548 443634 297600 443640
rect 297560 417081 297588 443634
rect 297652 421841 297680 443838
rect 298006 443592 298062 443601
rect 298006 443527 298062 443536
rect 298020 443018 298048 443527
rect 298008 443012 298060 443018
rect 298008 442954 298060 442960
rect 298008 431928 298060 431934
rect 298008 431870 298060 431876
rect 298020 430681 298048 431870
rect 298006 430672 298062 430681
rect 298006 430607 298062 430616
rect 298008 426420 298060 426426
rect 298008 426362 298060 426368
rect 298020 425921 298048 426362
rect 298006 425912 298062 425921
rect 298006 425847 298062 425856
rect 297638 421832 297694 421841
rect 297638 421767 297694 421776
rect 297546 417072 297602 417081
rect 297546 417007 297602 417016
rect 297454 412992 297510 413001
rect 297454 412927 297510 412936
rect 297362 408232 297418 408241
rect 297362 408167 297418 408176
rect 298008 404320 298060 404326
rect 298008 404262 298060 404268
rect 298020 404161 298048 404262
rect 298006 404152 298062 404161
rect 298006 404087 298062 404096
rect 297180 401396 297232 401402
rect 297180 401338 297232 401344
rect 297192 400994 297220 401338
rect 298008 401124 298060 401130
rect 298008 401066 298060 401072
rect 297180 400988 297232 400994
rect 297180 400930 297232 400936
rect 298020 400722 298048 401066
rect 298008 400716 298060 400722
rect 298008 400658 298060 400664
rect 298572 400178 298600 446150
rect 298652 444576 298704 444582
rect 298652 444518 298704 444524
rect 298560 400172 298612 400178
rect 298560 400114 298612 400120
rect 298664 398342 298692 444518
rect 298742 443864 298798 443873
rect 298742 443799 298798 443808
rect 298652 398336 298704 398342
rect 298652 398278 298704 398284
rect 298100 389972 298152 389978
rect 298100 389914 298152 389920
rect 296628 325644 296680 325650
rect 296628 325586 296680 325592
rect 296536 313268 296588 313274
rect 296536 313210 296588 313216
rect 296444 273216 296496 273222
rect 296444 273158 296496 273164
rect 296352 259412 296404 259418
rect 296352 259354 296404 259360
rect 296260 219428 296312 219434
rect 296260 219370 296312 219376
rect 296168 179376 296220 179382
rect 296168 179318 296220 179324
rect 296076 100700 296128 100706
rect 296076 100642 296128 100648
rect 296720 18896 296772 18902
rect 296720 18838 296772 18844
rect 296732 16574 296760 18838
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 291396 480 291424 16546
rect 292578 6624 292634 6633
rect 292578 6559 292634 6568
rect 292592 480 292620 6559
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 296076 3800 296128 3806
rect 296076 3742 296128 3748
rect 296088 480 296116 3742
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 389914
rect 298756 33114 298784 443799
rect 298848 113150 298876 446247
rect 298926 443184 298982 443193
rect 298926 443119 298982 443128
rect 298940 153202 298968 443119
rect 299032 233238 299060 446286
rect 299110 443320 299166 443329
rect 299110 443255 299166 443264
rect 299124 245614 299152 443255
rect 299216 379506 299244 447102
rect 299294 443456 299350 443465
rect 299294 443391 299350 443400
rect 299204 379500 299256 379506
rect 299204 379442 299256 379448
rect 299308 353258 299336 443391
rect 299400 398750 299428 448559
rect 299860 446486 299888 453478
rect 299848 446480 299900 446486
rect 299848 446422 299900 446428
rect 299480 445052 299532 445058
rect 299480 444994 299532 445000
rect 299492 422294 299520 444994
rect 299848 444440 299900 444446
rect 299848 444382 299900 444388
rect 299492 422266 299796 422294
rect 299664 400784 299716 400790
rect 299664 400726 299716 400732
rect 299388 398744 299440 398750
rect 299388 398686 299440 398692
rect 299676 398410 299704 400726
rect 299768 400466 299796 422266
rect 299860 400790 299888 444382
rect 383856 431954 383884 454022
rect 383934 453999 383990 454008
rect 384040 452305 384068 455534
rect 384026 452296 384082 452305
rect 384026 452231 384082 452240
rect 384132 452146 384160 455738
rect 384212 455728 384264 455734
rect 384212 455670 384264 455676
rect 383948 452118 384160 452146
rect 383948 438705 383976 452118
rect 384224 451274 384252 455670
rect 385040 455660 385092 455666
rect 385040 455602 385092 455608
rect 384304 455524 384356 455530
rect 384304 455466 384356 455472
rect 384040 451246 384252 451274
rect 384040 448225 384068 451246
rect 384026 448216 384082 448225
rect 384026 448151 384082 448160
rect 383934 438696 383990 438705
rect 383934 438631 383990 438640
rect 383856 431926 383976 431954
rect 384316 431934 384344 455466
rect 383948 421705 383976 431926
rect 384304 431928 384356 431934
rect 384304 431870 384356 431876
rect 383934 421696 383990 421705
rect 383934 421631 383990 421640
rect 385052 416401 385080 455602
rect 385144 430001 385172 455874
rect 385224 455864 385276 455870
rect 385224 455806 385276 455812
rect 385236 434081 385264 455806
rect 385328 442921 385356 456826
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580264 455456 580316 455462
rect 580264 455398 580316 455404
rect 385314 442912 385370 442921
rect 385314 442847 385370 442856
rect 385222 434072 385278 434081
rect 385222 434007 385278 434016
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 385130 429992 385186 430001
rect 385130 429927 385186 429936
rect 580276 418305 580304 455398
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 385038 416392 385094 416401
rect 385038 416327 385094 416336
rect 385038 407552 385094 407561
rect 385038 407487 385094 407496
rect 385052 401606 385080 407487
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 385040 401600 385092 401606
rect 385040 401542 385092 401548
rect 299848 400784 299900 400790
rect 382738 400752 382794 400761
rect 299848 400726 299900 400732
rect 307588 400722 307786 400738
rect 324240 400722 324530 400738
rect 332520 400722 332902 400738
rect 340984 400722 341274 400738
rect 307576 400716 307786 400722
rect 307628 400710 307786 400716
rect 324228 400716 324530 400722
rect 307576 400658 307628 400664
rect 324280 400710 324530 400716
rect 332508 400716 332902 400722
rect 324228 400658 324280 400664
rect 332560 400710 332902 400716
rect 340972 400716 341274 400722
rect 332508 400658 332560 400664
rect 341024 400710 341274 400716
rect 382794 400710 383134 400738
rect 382738 400687 382794 400696
rect 340972 400658 341024 400664
rect 299768 400438 300058 400466
rect 390558 400344 390614 400353
rect 390558 400279 390614 400288
rect 303908 398818 303936 400044
rect 303896 398812 303948 398818
rect 303896 398754 303948 398760
rect 299664 398404 299716 398410
rect 299664 398346 299716 398352
rect 312280 398274 312308 400044
rect 316144 398585 316172 400044
rect 316130 398576 316186 398585
rect 316130 398511 316186 398520
rect 320652 398342 320680 400044
rect 329024 399129 329052 400044
rect 329010 399120 329066 399129
rect 329010 399055 329066 399064
rect 337396 398857 337424 400044
rect 337382 398848 337438 398857
rect 337382 398783 337438 398792
rect 345768 398410 345796 400044
rect 349632 398478 349660 400044
rect 354140 398546 354168 400044
rect 358004 398614 358032 400044
rect 362512 398682 362540 400044
rect 362500 398676 362552 398682
rect 362500 398618 362552 398624
rect 357992 398608 358044 398614
rect 357992 398550 358044 398556
rect 354128 398540 354180 398546
rect 354128 398482 354180 398488
rect 349620 398472 349672 398478
rect 349620 398414 349672 398420
rect 345756 398404 345808 398410
rect 345756 398346 345808 398352
rect 320640 398336 320692 398342
rect 320640 398278 320692 398284
rect 312268 398268 312320 398274
rect 312268 398210 312320 398216
rect 366376 398206 366404 400044
rect 370884 398750 370912 400044
rect 370872 398744 370924 398750
rect 374748 398721 374776 400044
rect 370872 398686 370924 398692
rect 374734 398712 374790 398721
rect 374734 398647 374790 398656
rect 366364 398200 366416 398206
rect 366364 398142 366416 398148
rect 379256 397905 379284 400044
rect 379242 397896 379298 397905
rect 379242 397831 379298 397840
rect 310518 397352 310574 397361
rect 310518 397287 310574 397296
rect 305000 394528 305052 394534
rect 305000 394470 305052 394476
rect 299296 353252 299348 353258
rect 299296 353194 299348 353200
rect 299112 245608 299164 245614
rect 299112 245550 299164 245556
rect 299020 233232 299072 233238
rect 299020 233174 299072 233180
rect 298928 153196 298980 153202
rect 298928 153138 298980 153144
rect 298836 113144 298888 113150
rect 298836 113086 298888 113092
rect 298744 33108 298796 33114
rect 298744 33050 298796 33056
rect 300860 25764 300912 25770
rect 300860 25706 300912 25712
rect 299572 18828 299624 18834
rect 299572 18770 299624 18776
rect 299584 3398 299612 18770
rect 300872 16574 300900 25706
rect 303620 18760 303672 18766
rect 303620 18702 303672 18708
rect 303632 16574 303660 18702
rect 305012 16574 305040 394470
rect 307758 25528 307814 25537
rect 307758 25463 307814 25472
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299664 3732 299716 3738
rect 299664 3674 299716 3680
rect 299572 3392 299624 3398
rect 299572 3334 299624 3340
rect 299676 480 299704 3674
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303158 4040 303214 4049
rect 303158 3975 303214 3984
rect 303172 480 303200 3975
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 7812 306800 7818
rect 306748 7754 306800 7760
rect 306760 480 306788 7754
rect 307772 3398 307800 25463
rect 307850 18592 307906 18601
rect 307850 18527 307906 18536
rect 307864 16574 307892 18527
rect 310532 16574 310560 397287
rect 324318 397216 324374 397225
rect 324318 397151 324374 397160
rect 322940 394460 322992 394466
rect 322940 394402 322992 394408
rect 316040 352708 316092 352714
rect 316040 352650 316092 352656
rect 311900 87780 311952 87786
rect 311900 87722 311952 87728
rect 311912 16574 311940 87722
rect 314660 18692 314712 18698
rect 314660 18634 314712 18640
rect 307864 16546 307984 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 16546
rect 310242 7712 310298 7721
rect 310242 7647 310298 7656
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 7647
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313830 3904 313886 3913
rect 313830 3839 313886 3848
rect 313844 480 313872 3839
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 18634
rect 316052 16574 316080 352650
rect 318800 25696 318852 25702
rect 318800 25638 318852 25644
rect 317420 20324 317472 20330
rect 317420 20266 317472 20272
rect 317432 16574 317460 20266
rect 318812 16574 318840 25638
rect 321560 20256 321612 20262
rect 321560 20198 321612 20204
rect 321572 16574 321600 20198
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 321572 16546 322152 16574
rect 316236 480 316264 16546
rect 317328 6724 317380 6730
rect 317328 6666 317380 6672
rect 317340 480 317368 6666
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 320916 7744 320968 7750
rect 320916 7686 320968 7692
rect 320928 480 320956 7686
rect 322124 480 322152 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 394402
rect 324332 3398 324360 397151
rect 364338 397080 364394 397089
rect 364338 397015 364394 397024
rect 342260 396976 342312 396982
rect 342260 396918 342312 396924
rect 329840 394392 329892 394398
rect 329840 394334 329892 394340
rect 328458 83464 328514 83473
rect 328458 83399 328514 83408
rect 328472 16574 328500 83399
rect 329852 16574 329880 394334
rect 332600 394324 332652 394330
rect 332600 394266 332652 394272
rect 331220 391604 331272 391610
rect 331220 391546 331272 391552
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 326802 9072 326858 9081
rect 326802 9007 326858 9016
rect 324412 7676 324464 7682
rect 324412 7618 324464 7624
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 7618
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 326816 480 326844 9007
rect 327998 7576 328054 7585
rect 327998 7511 328054 7520
rect 328012 480 328040 7511
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 391546
rect 332612 3398 332640 394266
rect 340880 394188 340932 394194
rect 340880 394130 340932 394136
rect 336740 25628 336792 25634
rect 336740 25570 336792 25576
rect 336752 16574 336780 25570
rect 340892 16574 340920 394130
rect 342272 16574 342300 396918
rect 347780 394256 347832 394262
rect 347780 394198 347832 394204
rect 343638 27024 343694 27033
rect 343638 26959 343694 26968
rect 343652 16574 343680 26959
rect 346398 19952 346454 19961
rect 346398 19887 346454 19896
rect 346412 16574 346440 19887
rect 347792 16574 347820 394198
rect 357440 354272 357492 354278
rect 357440 354214 357492 354220
rect 353300 177472 353352 177478
rect 353300 177414 353352 177420
rect 350540 27260 350592 27266
rect 350540 27202 350592 27208
rect 349160 20188 349212 20194
rect 349160 20130 349212 20136
rect 336752 16546 337056 16574
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 332692 6656 332744 6662
rect 332692 6598 332744 6604
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 6598
rect 336280 6588 336332 6594
rect 336280 6530 336332 6536
rect 335084 3664 335136 3670
rect 335084 3606 335136 3612
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 3606
rect 336292 480 336320 6530
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 339866 6352 339922 6361
rect 339866 6287 339922 6296
rect 338670 3768 338726 3777
rect 338670 3703 338726 3712
rect 338684 480 338712 3703
rect 339880 480 339908 6287
rect 340984 480 341012 16546
rect 342168 6520 342220 6526
rect 342168 6462 342220 6468
rect 342180 480 342208 6462
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 345754 6488 345810 6497
rect 345754 6423 345810 6432
rect 345768 480 345796 6423
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3398 349200 20130
rect 350552 16574 350580 27202
rect 353312 16574 353340 177414
rect 354680 27192 354732 27198
rect 354680 27134 354732 27140
rect 354692 16574 354720 27134
rect 350552 16546 351224 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 349252 9308 349304 9314
rect 349252 9250 349304 9256
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 9250
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352840 9240 352892 9246
rect 352840 9182 352892 9188
rect 352852 480 352880 9182
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356336 9172 356388 9178
rect 356336 9114 356388 9120
rect 356348 480 356376 9114
rect 357452 3398 357480 354214
rect 360198 352880 360254 352889
rect 360198 352815 360254 352824
rect 357532 351280 357584 351286
rect 357532 351222 357584 351228
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 351222
rect 360212 16574 360240 352815
rect 361578 26888 361634 26897
rect 361578 26823 361634 26832
rect 361592 16574 361620 26823
rect 364352 16574 364380 397015
rect 372620 394120 372672 394126
rect 372620 394062 372672 394068
rect 365720 391536 365772 391542
rect 365720 391478 365772 391484
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 364352 16546 364656 16574
rect 359924 9104 359976 9110
rect 359924 9046 359976 9052
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 359936 480 359964 9046
rect 361132 480 361160 16546
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363510 8936 363566 8945
rect 363510 8871 363566 8880
rect 363524 480 363552 8871
rect 364628 480 364656 16546
rect 365732 1154 365760 391478
rect 365812 82272 365864 82278
rect 365812 82214 365864 82220
rect 365720 1148 365772 1154
rect 365720 1090 365772 1096
rect 365824 480 365852 82214
rect 368480 27124 368532 27130
rect 368480 27066 368532 27072
rect 367100 20120 367152 20126
rect 367100 20062 367152 20068
rect 367112 16574 367140 20062
rect 368492 16574 368520 27066
rect 371240 20052 371292 20058
rect 371240 19994 371292 20000
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 367008 1148 367060 1154
rect 367008 1090 367060 1096
rect 367020 480 367048 1090
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370596 9036 370648 9042
rect 370596 8978 370648 8984
rect 370608 480 370636 8978
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 19994
rect 372632 16574 372660 394062
rect 382280 394052 382332 394058
rect 382280 393994 382332 394000
rect 375380 87712 375432 87718
rect 375380 87654 375432 87660
rect 374000 19984 374052 19990
rect 374000 19926 374052 19932
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3398 374040 19926
rect 375392 16574 375420 87654
rect 378138 21720 378194 21729
rect 378138 21655 378194 21664
rect 378152 16574 378180 21655
rect 375392 16546 376064 16574
rect 378152 16546 378456 16574
rect 374092 10668 374144 10674
rect 374092 10610 374144 10616
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 10610
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377680 10464 377732 10470
rect 377680 10406 377732 10412
rect 377692 480 377720 10406
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 381174 10568 381230 10577
rect 379520 10532 379572 10538
rect 381174 10503 381230 10512
rect 379520 10474 379572 10480
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 10474
rect 381188 480 381216 10503
rect 382292 3398 382320 393994
rect 387800 391468 387852 391474
rect 387800 391410 387852 391416
rect 385040 352640 385092 352646
rect 385040 352582 385092 352588
rect 382370 21584 382426 21593
rect 382370 21519 382426 21528
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 21519
rect 385052 16574 385080 352582
rect 386420 27056 386472 27062
rect 386420 26998 386472 27004
rect 386432 16574 386460 26998
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 384304 10600 384356 10606
rect 384304 10542 384356 10548
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 10542
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 391410
rect 389180 17468 389232 17474
rect 389180 17410 389232 17416
rect 389192 16574 389220 17410
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 1154 390600 400279
rect 580000 400178 580028 404903
rect 579988 400172 580040 400178
rect 579988 400114 580040 400120
rect 437480 399016 437532 399022
rect 437480 398958 437532 398964
rect 398838 396944 398894 396953
rect 398838 396879 398894 396888
rect 402980 396908 403032 396914
rect 391940 389904 391992 389910
rect 391940 389846 391992 389852
rect 391952 16574 391980 389846
rect 393320 354204 393372 354210
rect 393320 354146 393372 354152
rect 393332 16574 393360 354146
rect 394700 177404 394752 177410
rect 394700 177346 394752 177352
rect 394712 16574 394740 177346
rect 397460 26988 397512 26994
rect 397460 26930 397512 26936
rect 396080 21684 396132 21690
rect 396080 21626 396132 21632
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390652 12164 390704 12170
rect 390652 12106 390704 12112
rect 390560 1148 390612 1154
rect 390560 1090 390612 1096
rect 390664 480 390692 12106
rect 391848 1148 391900 1154
rect 391848 1090 391900 1096
rect 391860 480 391888 1090
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 21626
rect 397472 16574 397500 26930
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3398 398880 396879
rect 402980 396850 403032 396856
rect 401600 392692 401652 392698
rect 401600 392634 401652 392640
rect 398930 351112 398986 351121
rect 398930 351047 398986 351056
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 351047
rect 400220 60104 400272 60110
rect 400220 60046 400272 60052
rect 400232 16574 400260 60046
rect 401612 16574 401640 392634
rect 402992 16574 403020 396850
rect 409880 396840 409932 396846
rect 409880 396782 409932 396788
rect 431958 396808 432014 396817
rect 407120 60036 407172 60042
rect 407120 59978 407172 59984
rect 404360 26920 404412 26926
rect 404360 26862 404412 26868
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 26862
rect 406016 10396 406068 10402
rect 406016 10338 406068 10344
rect 406028 480 406056 10338
rect 407132 3398 407160 59978
rect 407212 21616 407264 21622
rect 407212 21558 407264 21564
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 21558
rect 409892 16574 409920 396782
rect 431958 396743 432014 396752
rect 423680 352572 423732 352578
rect 423680 352514 423732 352520
rect 411260 87644 411312 87650
rect 411260 87586 411312 87592
rect 411272 16574 411300 87586
rect 420920 82204 420972 82210
rect 420920 82146 420972 82152
rect 414018 21448 414074 21457
rect 414018 21383 414074 21392
rect 414032 16574 414060 21383
rect 416778 21312 416834 21321
rect 416778 21247 416834 21256
rect 416792 16574 416820 21247
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 414032 16546 414336 16574
rect 416792 16546 417464 16574
rect 409144 10328 409196 10334
rect 409144 10270 409196 10276
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 10270
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 412638 10432 412694 10441
rect 412638 10367 412694 10376
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 10367
rect 414308 480 414336 16546
rect 415398 10296 415454 10305
rect 415398 10231 415454 10240
rect 415412 3398 415440 10231
rect 415492 8968 415544 8974
rect 415492 8910 415544 8916
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 8910
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418988 6452 419040 6458
rect 418988 6394 419040 6400
rect 419000 480 419028 6394
rect 420184 6384 420236 6390
rect 420184 6326 420236 6332
rect 420196 480 420224 6326
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 82146
rect 422576 14952 422628 14958
rect 422576 14894 422628 14900
rect 422588 480 422616 14894
rect 423692 1426 423720 352514
rect 429200 304292 429252 304298
rect 429200 304234 429252 304240
rect 427820 86556 427872 86562
rect 427820 86498 427872 86504
rect 427832 16574 427860 86498
rect 427832 16546 428504 16574
rect 425704 13524 425756 13530
rect 425704 13466 425756 13472
rect 423772 12096 423824 12102
rect 423772 12038 423824 12044
rect 423680 1420 423732 1426
rect 423680 1362 423732 1368
rect 423784 480 423812 12038
rect 424968 1420 425020 1426
rect 424968 1362 425020 1368
rect 424980 480 425008 1362
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 13466
rect 426808 12028 426860 12034
rect 426808 11970 426860 11976
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 11970
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 304234
rect 430856 11960 430908 11966
rect 430856 11902 430908 11908
rect 430868 480 430896 11902
rect 431972 1170 432000 396743
rect 436100 333260 436152 333266
rect 436100 333202 436152 333208
rect 434718 177304 434774 177313
rect 434718 177239 434774 177248
rect 434732 16574 434760 177239
rect 436112 16574 436140 333202
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432050 16280 432106 16289
rect 432050 16215 432106 16224
rect 432064 3398 432092 16215
rect 433982 11792 434038 11801
rect 433982 11727 434038 11736
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 11727
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 398958
rect 543740 398948 543792 398954
rect 543740 398890 543792 398896
rect 489918 398304 489974 398313
rect 489918 398239 489974 398248
rect 480260 398132 480312 398138
rect 480260 398074 480312 398080
rect 473360 396772 473412 396778
rect 473360 396714 473412 396720
rect 452658 396672 452714 396681
rect 452658 396607 452714 396616
rect 440240 391400 440292 391406
rect 440240 391342 440292 391348
rect 438860 21548 438912 21554
rect 438860 21490 438912 21496
rect 438872 16574 438900 21490
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 391342
rect 445760 355428 445812 355434
rect 445760 355370 445812 355376
rect 440332 354136 440384 354142
rect 440332 354078 440384 354084
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 354078
rect 443000 180124 443052 180130
rect 443000 180066 443052 180072
rect 441620 21480 441672 21486
rect 441620 21422 441672 21428
rect 441632 16574 441660 21422
rect 443012 16574 443040 180066
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445024 11892 445076 11898
rect 445024 11834 445076 11840
rect 445036 480 445064 11834
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 355370
rect 449900 182844 449952 182850
rect 449900 182786 449952 182792
rect 447140 86488 447192 86494
rect 447140 86430 447192 86436
rect 447152 16574 447180 86430
rect 448520 21412 448572 21418
rect 448520 21354 448572 21360
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 1426 448560 21354
rect 449912 16574 449940 182786
rect 452672 16574 452700 396607
rect 456800 391332 456852 391338
rect 456800 391274 456852 391280
rect 454040 86420 454092 86426
rect 454040 86362 454092 86368
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 448612 11824 448664 11830
rect 448612 11766 448664 11772
rect 448520 1420 448572 1426
rect 448520 1362 448572 1368
rect 448624 480 448652 11766
rect 449808 1420 449860 1426
rect 449808 1362 449860 1368
rect 449820 480 449848 1362
rect 450924 480 450952 16546
rect 451646 11656 451702 11665
rect 451646 11591 451702 11600
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 11591
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 86362
rect 455696 11756 455748 11762
rect 455696 11698 455748 11704
rect 455708 480 455736 11698
rect 456812 3210 456840 391274
rect 470598 82104 470654 82113
rect 470598 82039 470654 82048
rect 467840 31068 467892 31074
rect 467840 31010 467892 31016
rect 460940 29640 460992 29646
rect 460940 29582 460992 29588
rect 456892 28280 456944 28286
rect 456892 28222 456944 28228
rect 456904 3398 456932 28222
rect 459560 23180 459612 23186
rect 459560 23122 459612 23128
rect 459572 16574 459600 23122
rect 460952 16574 460980 29582
rect 463700 23112 463752 23118
rect 463700 23054 463752 23060
rect 463712 16574 463740 23054
rect 466458 22808 466514 22817
rect 466458 22743 466514 22752
rect 466472 16574 466500 22743
rect 467852 16574 467880 31010
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 459192 13456 459244 13462
rect 459192 13398 459244 13404
rect 456892 3392 456944 3398
rect 456892 3334 456944 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 456812 3182 456932 3210
rect 456904 480 456932 3182
rect 458100 480 458128 3334
rect 459204 480 459232 13398
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 462320 13388 462372 13394
rect 462320 13330 462372 13336
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 13330
rect 463988 480 464016 16546
rect 465816 13320 465868 13326
rect 465816 13262 465868 13268
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 465184 480 465212 3538
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 13262
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469862 13152 469918 13161
rect 469862 13087 469918 13096
rect 469876 480 469904 13087
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 82039
rect 471980 18624 472032 18630
rect 471980 18566 472032 18572
rect 471992 16574 472020 18566
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3602 473400 396714
rect 474740 184204 474792 184210
rect 474740 184146 474792 184152
rect 474752 16574 474780 184146
rect 478880 86352 478932 86358
rect 478880 86294 478932 86300
rect 477500 23044 477552 23050
rect 477500 22986 477552 22992
rect 477512 16574 477540 22986
rect 474752 16546 475792 16574
rect 477512 16546 478184 16574
rect 473452 13252 473504 13258
rect 473452 13194 473504 13200
rect 473360 3596 473412 3602
rect 473360 3538 473412 3544
rect 473464 480 473492 13194
rect 474188 3596 474240 3602
rect 474188 3538 474240 3544
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3538
rect 475764 480 475792 16546
rect 476488 13184 476540 13190
rect 476488 13126 476540 13132
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 13126
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 86294
rect 480272 16574 480300 398074
rect 483018 397488 483074 397497
rect 483018 397423 483074 397432
rect 481640 22976 481692 22982
rect 481640 22918 481692 22924
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 3602 481680 22918
rect 483032 16574 483060 397423
rect 488538 354240 488594 354249
rect 488538 354175 488594 354184
rect 485778 22672 485834 22681
rect 485778 22607 485834 22616
rect 485792 16574 485820 22607
rect 488552 16574 488580 354175
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 481732 13116 481784 13122
rect 481732 13058 481784 13064
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 13058
rect 482468 3596 482520 3602
rect 482468 3538 482520 3544
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3538
rect 484044 480 484072 16546
rect 484766 13016 484822 13025
rect 484766 12951 484822 12960
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 12951
rect 486436 480 486464 16546
rect 487618 3632 487674 3641
rect 487618 3567 487674 3576
rect 487632 480 487660 3567
rect 488828 480 488856 16546
rect 489932 3602 489960 398239
rect 494058 398168 494114 398177
rect 494058 398103 494114 398112
rect 490012 22908 490064 22914
rect 490012 22850 490064 22856
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 490024 3482 490052 22850
rect 492680 22840 492732 22846
rect 492680 22782 492732 22788
rect 492692 16574 492720 22782
rect 494072 16574 494100 398103
rect 507858 398032 507914 398041
rect 507858 397967 507914 397976
rect 498200 392624 498252 392630
rect 498200 392566 498252 392572
rect 496820 177336 496872 177342
rect 496820 177278 496872 177284
rect 496832 16574 496860 177278
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 492312 14884 492364 14890
rect 492312 14826 492364 14832
rect 490748 3596 490800 3602
rect 490748 3538 490800 3544
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3538
rect 492324 480 492352 14826
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 495440 14816 495492 14822
rect 495440 14758 495492 14764
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 14758
rect 497108 480 497136 16546
rect 498212 480 498240 392566
rect 499580 389836 499632 389842
rect 499580 389778 499632 389784
rect 499592 16574 499620 389778
rect 506478 352744 506534 352753
rect 506478 352679 506534 352688
rect 503718 24304 503774 24313
rect 503718 24239 503774 24248
rect 499592 16546 500632 16574
rect 498936 14748 498988 14754
rect 498936 14690 498988 14696
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 14690
rect 500604 480 500632 16546
rect 502984 14680 503036 14686
rect 502984 14622 503036 14628
rect 501788 3528 501840 3534
rect 501788 3470 501840 3476
rect 501800 480 501828 3470
rect 502996 480 503024 14622
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 24239
rect 505374 3496 505430 3505
rect 505374 3431 505430 3440
rect 505388 480 505416 3431
rect 506492 480 506520 352679
rect 506572 22772 506624 22778
rect 506572 22714 506624 22720
rect 506584 16574 506612 22714
rect 507872 16574 507900 397967
rect 525800 397520 525852 397526
rect 525800 397462 525852 397468
rect 521658 395448 521714 395457
rect 521658 395383 521714 395392
rect 512000 391264 512052 391270
rect 512000 391206 512052 391212
rect 510620 24472 510672 24478
rect 510620 24414 510672 24420
rect 510632 16574 510660 24414
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 509608 14612 509660 14618
rect 509608 14554 509660 14560
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 14554
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 391206
rect 514760 355360 514812 355366
rect 514760 355302 514812 355308
rect 513380 14544 513432 14550
rect 513380 14486 513432 14492
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 14486
rect 514772 3534 514800 355302
rect 517520 86284 517572 86290
rect 517520 86226 517572 86232
rect 514852 24404 514904 24410
rect 514852 24346 514904 24352
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 24346
rect 517532 16574 517560 86226
rect 517532 16546 517928 16574
rect 517152 14476 517204 14482
rect 517152 14418 517204 14424
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 14418
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 520278 14512 520334 14521
rect 520278 14447 520334 14456
rect 519544 5228 519596 5234
rect 519544 5170 519596 5176
rect 519556 480 519584 5170
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 14447
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 395383
rect 524420 24336 524472 24342
rect 524420 24278 524472 24284
rect 524432 16574 524460 24278
rect 525812 16574 525840 397462
rect 535460 395548 535512 395554
rect 535460 395490 535512 395496
rect 534080 354068 534132 354074
rect 534080 354010 534132 354016
rect 528560 24268 528612 24274
rect 528560 24210 528612 24216
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523774 16144 523830 16153
rect 523774 16079 523830 16088
rect 523038 4992 523094 5001
rect 523038 4927 523094 4936
rect 523052 480 523080 4927
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16079
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 16176 527876 16182
rect 527824 16118 527876 16124
rect 527836 480 527864 16118
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 24210
rect 531320 24200 531372 24206
rect 531320 24142 531372 24148
rect 531332 3534 531360 24142
rect 534092 16574 534120 354010
rect 535472 16574 535500 395490
rect 542360 395480 542412 395486
rect 542360 395422 542412 395428
rect 538218 354104 538274 354113
rect 538218 354039 538274 354048
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 531412 16108 531464 16114
rect 531412 16050 531464 16056
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 530124 3460 530176 3466
rect 530124 3402 530176 3408
rect 530136 480 530164 3402
rect 531424 3346 531452 16050
rect 533712 5160 533764 5166
rect 533712 5102 533764 5108
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 5102
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 5092 537260 5098
rect 537208 5034 537260 5040
rect 537220 480 537248 5034
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 354039
rect 539598 86184 539654 86193
rect 539598 86119 539654 86128
rect 539612 480 539640 86119
rect 542372 16574 542400 395422
rect 543752 16574 543780 398890
rect 564440 398880 564492 398886
rect 564440 398822 564492 398828
rect 549260 395412 549312 395418
rect 549260 395354 549312 395360
rect 546500 354000 546552 354006
rect 546500 353942 546552 353948
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 541990 16008 542046 16017
rect 541990 15943 542046 15952
rect 540794 4856 540850 4865
rect 540794 4791 540850 4800
rect 540808 480 540836 4791
rect 542004 480 542032 15943
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 16040 545540 16046
rect 545488 15982 545540 15988
rect 545500 480 545528 15982
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 353942
rect 549272 16574 549300 395354
rect 556158 395312 556214 395321
rect 556158 395247 556214 395256
rect 549272 16546 550312 16574
rect 548616 15972 548668 15978
rect 548616 15914 548668 15920
rect 547880 5024 547932 5030
rect 547880 4966 547932 4972
rect 547892 480 547920 4966
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 15914
rect 550284 480 550312 16546
rect 552664 15904 552716 15910
rect 552664 15846 552716 15852
rect 551468 4956 551520 4962
rect 551468 4898 551520 4904
rect 551480 480 551508 4898
rect 552676 480 552704 15846
rect 553768 7608 553820 7614
rect 553768 7550 553820 7556
rect 553780 480 553808 7550
rect 554964 4888 555016 4894
rect 554964 4830 555016 4836
rect 554976 480 555004 4830
rect 556172 3534 556200 395247
rect 557538 355328 557594 355337
rect 557538 355263 557594 355272
rect 557552 16574 557580 355263
rect 558918 353968 558974 353977
rect 558918 353903 558974 353912
rect 558932 16574 558960 353903
rect 563060 17400 563112 17406
rect 563060 17342 563112 17348
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 556250 15872 556306 15881
rect 556250 15807 556306 15816
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 15807
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 562048 6316 562100 6322
rect 562048 6258 562100 6264
rect 560852 4820 560904 4826
rect 560852 4762 560904 4768
rect 560864 480 560892 4762
rect 562060 480 562088 6258
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 17342
rect 564452 3534 564480 398822
rect 564532 395344 564584 395350
rect 564532 395286 564584 395292
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 395286
rect 571340 393984 571392 393990
rect 571340 393926 571392 393932
rect 567200 24132 567252 24138
rect 567200 24074 567252 24080
rect 565820 17332 565872 17338
rect 565820 17274 565872 17280
rect 565832 16574 565860 17274
rect 567212 16574 567240 24074
rect 569960 17264 570012 17270
rect 569960 17206 570012 17212
rect 569972 16574 570000 17206
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 6248 569184 6254
rect 569132 6190 569184 6196
rect 569144 480 569172 6190
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 393926
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 576858 352608 576914 352617
rect 576858 352543 576914 352552
rect 572720 351212 572772 351218
rect 572720 351154 572772 351160
rect 572732 16574 572760 351154
rect 574098 24168 574154 24177
rect 574098 24103 574154 24112
rect 574112 16574 574140 24103
rect 576872 16574 576900 352543
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 581000 334620 581052 334626
rect 581000 334562 581052 334568
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 578240 25560 578292 25566
rect 578240 25502 578292 25508
rect 578252 16574 578280 25502
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 572720 6180 572772 6186
rect 572720 6122 572772 6128
rect 572732 480 572760 6122
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576306 6216 576362 6225
rect 576306 6151 576362 6160
rect 576320 480 576348 6151
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 581012 3534 581040 334562
rect 582380 185632 582432 185638
rect 582380 185574 582432 185580
rect 581092 82136 581144 82142
rect 581092 82078 581144 82084
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 579802 3360 579858 3369
rect 581104 3346 581132 82078
rect 582392 16574 582420 185574
rect 582392 16546 583432 16574
rect 581828 3528 581880 3534
rect 581828 3470 581880 3476
rect 579802 3295 579858 3304
rect 581012 3318 581132 3346
rect 579816 480 579844 3295
rect 581012 480 581040 3318
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581840 354 581868 3470
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581840 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 566888 3386 566944
rect 3146 553832 3202 553888
rect 3330 527856 3386 527912
rect 3238 501744 3294 501800
rect 3238 475632 3294 475688
rect 2870 462576 2926 462632
rect 3238 449520 3294 449576
rect 3514 671200 3570 671256
rect 3606 658144 3662 658200
rect 3698 632032 3754 632088
rect 3790 619112 3846 619168
rect 3882 606056 3938 606112
rect 3974 579944 4030 580000
rect 4066 514800 4122 514856
rect 78586 636384 78642 636440
rect 78310 635296 78366 635352
rect 78218 633664 78274 633720
rect 77758 632576 77814 632632
rect 78126 630944 78182 631000
rect 77850 629584 77906 629640
rect 77758 523504 77814 523560
rect 77666 520920 77722 520976
rect 78034 627952 78090 628008
rect 77942 608640 77998 608696
rect 77850 521600 77906 521656
rect 78402 610000 78458 610056
rect 78494 607688 78550 607744
rect 102874 597488 102930 597544
rect 111706 597488 111762 597544
rect 92478 597352 92534 597408
rect 100666 597352 100722 597408
rect 99286 597216 99342 597272
rect 94042 597080 94098 597136
rect 104806 597236 104862 597272
rect 104806 597216 104808 597236
rect 104808 597216 104860 597236
rect 104860 597216 104862 597236
rect 78494 526632 78550 526688
rect 78310 526496 78366 526552
rect 78310 523640 78366 523696
rect 78126 521600 78182 521656
rect 78126 520240 78182 520296
rect 78034 499840 78090 499896
rect 77942 498616 77998 498672
rect 78402 498344 78458 498400
rect 78586 517928 78642 517984
rect 102046 597080 102102 597136
rect 103426 596944 103482 597000
rect 106186 596964 106242 597000
rect 106186 596944 106188 596964
rect 106188 596944 106240 596964
rect 106240 596944 106242 596964
rect 97906 596828 97962 596864
rect 97906 596808 97908 596828
rect 97908 596808 97960 596828
rect 97960 596808 97962 596828
rect 95238 596264 95294 596320
rect 131026 596944 131082 597000
rect 126886 596672 126942 596728
rect 136546 596536 136602 596592
rect 140686 596556 140742 596592
rect 140686 596536 140688 596556
rect 140688 596536 140740 596556
rect 140740 596536 140742 596556
rect 115846 596264 115902 596320
rect 121366 596284 121422 596320
rect 121366 596264 121368 596284
rect 121368 596264 121420 596284
rect 121420 596264 121422 596284
rect 92938 488452 92940 488472
rect 92940 488452 92992 488472
rect 92992 488452 92994 488472
rect 92938 488416 92994 488452
rect 94226 488436 94282 488472
rect 94226 488416 94228 488436
rect 94228 488416 94280 488436
rect 94280 488416 94282 488436
rect 95330 488416 95386 488472
rect 97814 488416 97870 488472
rect 98918 488416 98974 488472
rect 100022 488416 100078 488472
rect 101126 488416 101182 488472
rect 102414 488416 102470 488472
rect 104806 488416 104862 488472
rect 105726 488416 105782 488472
rect 105818 488144 105874 488200
rect 111706 488144 111762 488200
rect 103426 487892 103482 487928
rect 103426 487872 103428 487892
rect 103428 487872 103480 487892
rect 103480 487872 103482 487892
rect 115846 487192 115902 487248
rect 121366 487192 121422 487248
rect 126886 487192 126942 487248
rect 131026 487192 131082 487248
rect 136546 487192 136602 487248
rect 140686 487192 140742 487248
rect 173162 596808 173218 596864
rect 187330 637064 187386 637120
rect 186778 635976 186834 636032
rect 186870 634344 186926 634400
rect 187238 631624 187294 631680
rect 187146 628632 187202 628688
rect 187054 610272 187110 610328
rect 186962 608368 187018 608424
rect 186778 525952 186834 526008
rect 186870 524320 186926 524376
rect 186778 523232 186834 523288
rect 186686 498208 186742 498264
rect 186870 521464 186926 521520
rect 186870 520240 186926 520296
rect 187422 633256 187478 633312
rect 187330 527040 187386 527096
rect 187330 524320 187386 524376
rect 187238 521600 187294 521656
rect 187146 518608 187202 518664
rect 187054 500248 187110 500304
rect 186962 498208 187018 498264
rect 187514 630264 187570 630320
rect 187422 523232 187478 523288
rect 187606 608640 187662 608696
rect 187514 521464 187570 521520
rect 187606 498616 187662 498672
rect 188434 525952 188490 526008
rect 3238 423544 3294 423600
rect 2778 410488 2834 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3146 267144 3202 267200
rect 3054 214920 3110 214976
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3146 110608 3202 110664
rect 2778 97552 2834 97608
rect 3514 446392 3570 446448
rect 3422 84632 3478 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 4066 345344 4122 345400
rect 3974 254088 4030 254144
rect 3882 241032 3938 241088
rect 3790 201864 3846 201920
rect 3698 188808 3754 188864
rect 3606 136720 3662 136776
rect 3514 45464 3570 45520
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 207846 597488 207902 597544
rect 208950 597488 209006 597544
rect 209962 597488 210018 597544
rect 211158 597488 211214 597544
rect 212354 597488 212410 597544
rect 213826 597488 213882 597544
rect 214838 597488 214894 597544
rect 215298 597488 215354 597544
rect 215758 597488 215814 597544
rect 226246 597488 226302 597544
rect 235906 597488 235962 597544
rect 245566 597488 245622 597544
rect 251086 597488 251142 597544
rect 204350 597080 204406 597136
rect 202878 596400 202934 596456
rect 204258 596264 204314 596320
rect 219438 596264 219494 596320
rect 189078 498616 189134 498672
rect 231766 597216 231822 597272
rect 241426 596808 241482 596864
rect 204718 488436 204774 488472
rect 204718 488416 204720 488436
rect 204720 488416 204772 488436
rect 204772 488416 204774 488436
rect 214838 488416 214894 488472
rect 202878 488180 202880 488200
rect 202880 488180 202932 488200
rect 202932 488180 202934 488200
rect 202878 488144 202934 488180
rect 211158 488280 211214 488336
rect 213734 488280 213790 488336
rect 203522 487192 203578 487248
rect 208858 487872 208914 487928
rect 215758 488280 215814 488336
rect 212354 487464 212410 487520
rect 204902 487192 204958 487248
rect 207662 487192 207718 487248
rect 210422 487212 210478 487248
rect 210422 487192 210424 487212
rect 210424 487192 210476 487212
rect 210476 487192 210478 487212
rect 216586 487192 216642 487248
rect 211158 447208 211214 447264
rect 210422 446256 210478 446312
rect 209134 446120 209190 446176
rect 79322 445984 79378 446040
rect 25502 397432 25558 397488
rect 13818 392536 13874 392592
rect 1674 9016 1730 9072
rect 570 8880 626 8936
rect 17038 11600 17094 11656
rect 27710 395256 27766 395312
rect 45558 395392 45614 395448
rect 30102 11736 30158 11792
rect 64878 396616 64934 396672
rect 63498 177248 63554 177304
rect 67638 395528 67694 395584
rect 50158 14456 50214 14512
rect 48502 11872 48558 11928
rect 51354 7520 51410 7576
rect 66718 12960 66774 13016
rect 188342 398248 188398 398304
rect 100758 396752 100814 396808
rect 84198 353912 84254 353968
rect 83278 10240 83334 10296
rect 86406 10376 86462 10432
rect 88246 9152 88302 9208
rect 88982 13096 89038 13152
rect 99838 15816 99894 15872
rect 118698 395664 118754 395720
rect 102138 354048 102194 354104
rect 120078 177384 120134 177440
rect 122286 12008 122342 12064
rect 139398 394032 139454 394088
rect 135258 393896 135314 393952
rect 138662 14592 138718 14648
rect 137650 7656 137706 7712
rect 138846 7792 138902 7848
rect 153198 394168 153254 394224
rect 151818 392672 151874 392728
rect 178682 398112 178738 398168
rect 173898 177520 173954 177576
rect 170310 15952 170366 16008
rect 173162 6160 173218 6216
rect 175462 3304 175518 3360
rect 187698 178608 187754 178664
rect 185582 10512 185638 10568
rect 191838 352552 191894 352608
rect 190458 46144 190514 46200
rect 194414 6296 194470 6352
rect 210054 444896 210110 444952
rect 209686 444760 209742 444816
rect 209502 444080 209558 444136
rect 209410 443808 209466 443864
rect 210238 444624 210294 444680
rect 210790 444488 210846 444544
rect 210606 444080 210662 444136
rect 209962 443536 210018 443592
rect 220726 487192 220782 487248
rect 226246 487192 226302 487248
rect 223302 446528 223358 446584
rect 224406 448568 224462 448624
rect 225694 454008 225750 454064
rect 225510 444080 225566 444136
rect 226246 445848 226302 445904
rect 226706 444080 226762 444136
rect 211066 443400 211122 443456
rect 212354 443400 212410 443456
rect 213642 443400 213698 443456
rect 226338 443672 226394 443728
rect 229742 446664 229798 446720
rect 229190 446392 229246 446448
rect 229374 445984 229430 446040
rect 231766 487192 231822 487248
rect 226706 443672 226762 443728
rect 231674 448704 231730 448760
rect 232042 454280 232098 454336
rect 232134 454144 232190 454200
rect 235906 487192 235962 487248
rect 241426 487192 241482 487248
rect 234066 449792 234122 449848
rect 238022 444080 238078 444136
rect 244646 487192 244702 487248
rect 249798 487192 249854 487248
rect 245474 443944 245530 444000
rect 250994 443944 251050 444000
rect 253478 444216 253534 444272
rect 254398 444352 254454 444408
rect 255410 449656 255466 449712
rect 255502 446392 255558 446448
rect 256422 449656 256478 449712
rect 293314 488416 293370 488472
rect 293866 488416 293922 488472
rect 293866 488008 293922 488064
rect 298006 636928 298062 636984
rect 297178 635840 297234 635896
rect 297086 610136 297142 610192
rect 296994 608640 297050 608696
rect 296902 517520 296958 517576
rect 297914 634208 297970 634264
rect 297730 633120 297786 633176
rect 297454 631488 297510 631544
rect 297178 525952 297234 526008
rect 297086 500248 297142 500304
rect 296902 488280 296958 488336
rect 292026 449656 292082 449712
rect 256422 444080 256478 444136
rect 256790 445712 256846 445768
rect 265622 444624 265678 444680
rect 203430 398792 203486 398848
rect 202142 398384 202198 398440
rect 203706 398656 203762 398712
rect 203522 398520 203578 398576
rect 203430 397432 203486 397488
rect 205822 398656 205878 398712
rect 205822 398384 205878 398440
rect 210330 397568 210386 397624
rect 210422 397432 210478 397488
rect 210422 397296 210478 397352
rect 209870 396344 209926 396400
rect 211158 398248 211214 398304
rect 211158 397840 211214 397896
rect 211250 397704 211306 397760
rect 211434 398248 211490 398304
rect 211342 397432 211398 397488
rect 211526 397976 211582 398032
rect 211618 397568 211674 397624
rect 211894 398656 211950 398712
rect 211802 398520 211858 398576
rect 211802 397568 211858 397624
rect 212446 397976 212502 398032
rect 212538 397704 212594 397760
rect 212630 397432 212686 397488
rect 212814 398384 212870 398440
rect 212998 397568 213054 397624
rect 213366 398112 213422 398168
rect 213918 399064 213974 399120
rect 214010 397976 214066 398032
rect 213918 397840 213974 397896
rect 214010 397568 214066 397624
rect 214286 397704 214342 397760
rect 214194 397568 214250 397624
rect 214102 397432 214158 397488
rect 214470 398928 214526 398984
rect 214470 398792 214526 398848
rect 215298 397432 215354 397488
rect 215574 397704 215630 397760
rect 215482 397568 215538 397624
rect 215390 396616 215446 396672
rect 215850 398112 215906 398168
rect 216678 397704 216734 397760
rect 216954 399200 217010 399256
rect 216862 397568 216918 397624
rect 216770 397432 216826 397488
rect 217046 397840 217102 397896
rect 218058 397432 218114 397488
rect 218242 397568 218298 397624
rect 218150 396752 218206 396808
rect 219530 397432 219586 397488
rect 219806 397568 219862 397624
rect 219714 397432 219770 397488
rect 219622 395664 219678 395720
rect 220910 397568 220966 397624
rect 221094 397568 221150 397624
rect 221002 397432 221058 397488
rect 221186 397432 221242 397488
rect 222198 397704 222254 397760
rect 222290 397432 222346 397488
rect 223578 397840 223634 397896
rect 223854 397704 223910 397760
rect 223946 397568 224002 397624
rect 223762 397432 223818 397488
rect 224958 397704 225014 397760
rect 225234 397568 225290 397624
rect 225142 397432 225198 397488
rect 225418 397840 225474 397896
rect 226430 396344 226486 396400
rect 229006 397840 229062 397896
rect 228914 397432 228970 397488
rect 230202 397976 230258 398032
rect 230386 397704 230442 397760
rect 230110 397568 230166 397624
rect 230018 397432 230074 397488
rect 231582 397704 231638 397760
rect 231766 397568 231822 397624
rect 231674 397432 231730 397488
rect 232962 397976 233018 398032
rect 232870 397568 232926 397624
rect 233146 397704 233202 397760
rect 233054 397432 233110 397488
rect 233882 398520 233938 398576
rect 234434 397704 234490 397760
rect 234342 397568 234398 397624
rect 234250 397432 234306 397488
rect 234526 397296 234582 397352
rect 234710 397840 234766 397896
rect 235722 397568 235778 397624
rect 235906 397704 235962 397760
rect 235814 397432 235870 397488
rect 235630 397160 235686 397216
rect 234894 5480 234950 5536
rect 236734 398112 236790 398168
rect 237102 397704 237158 397760
rect 237286 397568 237342 397624
rect 237194 397432 237250 397488
rect 237654 394440 237710 394496
rect 237838 394576 237894 394632
rect 238022 394440 238078 394496
rect 235998 3712 236054 3768
rect 237930 393896 237986 393952
rect 238390 397704 238446 397760
rect 238482 397568 238538 397624
rect 238574 397432 238630 397488
rect 238666 397024 238722 397080
rect 239218 394440 239274 394496
rect 239034 393896 239090 393952
rect 239770 397432 239826 397488
rect 240046 397568 240102 397624
rect 239954 397432 240010 397488
rect 240782 399880 240838 399936
rect 241334 397432 241390 397488
rect 241426 396888 241482 396944
rect 239310 3576 239366 3632
rect 240506 3440 240562 3496
rect 242530 397704 242586 397760
rect 242438 397568 242494 397624
rect 242806 397840 242862 397896
rect 242714 397432 242770 397488
rect 243910 398928 243966 398984
rect 244370 398656 244426 398712
rect 244186 397704 244242 397760
rect 244094 397568 244150 397624
rect 244002 397432 244058 397488
rect 244370 396752 244426 396808
rect 244186 393780 244242 393816
rect 244186 393760 244188 393780
rect 244188 393760 244240 393780
rect 244240 393760 244242 393780
rect 245474 397432 245530 397488
rect 245566 396616 245622 396672
rect 246210 393760 246266 393816
rect 246486 398248 246542 398304
rect 246670 397568 246726 397624
rect 246946 397704 247002 397760
rect 246854 397432 246910 397488
rect 247958 397976 248014 398032
rect 248142 397704 248198 397760
rect 248050 397568 248106 397624
rect 248326 397840 248382 397896
rect 248234 397432 248290 397488
rect 248510 399064 248566 399120
rect 248786 398520 248842 398576
rect 249522 397568 249578 397624
rect 249706 397704 249762 397760
rect 249614 397432 249670 397488
rect 249890 398112 249946 398168
rect 250166 398792 250222 398848
rect 250902 397840 250958 397896
rect 250810 397568 250866 397624
rect 251086 397704 251142 397760
rect 250810 397432 250866 397488
rect 250994 397432 251050 397488
rect 251270 398248 251326 398304
rect 252190 397840 252246 397896
rect 252282 397704 252338 397760
rect 252558 399200 252614 399256
rect 252466 397568 252522 397624
rect 252374 397432 252430 397488
rect 252650 398792 252706 398848
rect 252742 398656 252798 398712
rect 253202 397432 253258 397488
rect 253478 399880 253534 399936
rect 253570 397432 253626 397488
rect 253846 398384 253902 398440
rect 253754 397704 253810 397760
rect 254030 397976 254086 398032
rect 255042 397704 255098 397760
rect 255226 397840 255282 397896
rect 255134 397568 255190 397624
rect 254674 5072 254730 5128
rect 253478 3304 253534 3360
rect 256238 398248 256294 398304
rect 256054 397976 256110 398032
rect 255594 397840 255650 397896
rect 255318 395664 255374 395720
rect 257342 396480 257398 396536
rect 265806 443672 265862 443728
rect 273902 444896 273958 444952
rect 268382 444488 268438 444544
rect 273258 354320 273314 354376
rect 293130 442720 293186 442776
rect 292946 442448 293002 442504
rect 297546 628496 297602 628552
rect 297362 524320 297418 524376
rect 297638 608232 297694 608288
rect 297454 521600 297510 521656
rect 297546 518608 297602 518664
rect 297546 517520 297602 517576
rect 297822 630128 297878 630184
rect 317694 597488 317750 597544
rect 320086 597488 320142 597544
rect 320914 597488 320970 597544
rect 322202 597488 322258 597544
rect 322938 597488 322994 597544
rect 324318 597488 324374 597544
rect 326158 597488 326214 597544
rect 329838 597488 329894 597544
rect 345018 597488 345074 597544
rect 360198 597488 360254 597544
rect 313278 597216 313334 597272
rect 297822 524320 297878 524376
rect 297730 523232 297786 523288
rect 297638 498344 297694 498400
rect 297362 488416 297418 488472
rect 297362 488280 297418 488336
rect 298006 527040 298062 527096
rect 298006 520240 298062 520296
rect 297822 498616 297878 498672
rect 297914 489776 297970 489832
rect 297638 452376 297694 452432
rect 297822 488416 297878 488472
rect 297914 449792 297970 449848
rect 298006 448296 298062 448352
rect 295982 447208 296038 447264
rect 293130 400832 293186 400888
rect 293774 442584 293830 442640
rect 275282 397840 275338 397896
rect 291198 395528 291254 395584
rect 276018 6704 276074 6760
rect 274822 3168 274878 3224
rect 289818 18808 289874 18864
rect 292578 18672 292634 18728
rect 296074 442312 296130 442368
rect 314658 596828 314714 596864
rect 314658 596808 314660 596828
rect 314660 596808 314712 596828
rect 314712 596808 314714 596828
rect 319994 597352 320050 597408
rect 311898 596536 311954 596592
rect 324410 597352 324466 597408
rect 335358 597372 335414 597408
rect 335358 597352 335360 597372
rect 335360 597352 335412 597372
rect 335412 597352 335414 597372
rect 339498 596944 339554 597000
rect 349158 597080 349214 597136
rect 354678 596264 354734 596320
rect 314290 488416 314346 488472
rect 315394 488416 315450 488472
rect 313002 487872 313058 487928
rect 324410 487872 324466 487928
rect 319994 487484 320050 487520
rect 319994 487464 319996 487484
rect 319996 487464 320048 487484
rect 320048 487464 320050 487484
rect 322938 487464 322994 487520
rect 318062 487192 318118 487248
rect 319442 487192 319498 487248
rect 322202 487328 322258 487384
rect 320822 487212 320878 487248
rect 320822 487192 320824 487212
rect 320824 487192 320876 487212
rect 320876 487192 320878 487212
rect 326618 487736 326674 487792
rect 324318 487192 324374 487248
rect 329838 487192 329894 487248
rect 335358 487192 335414 487248
rect 339498 487192 339554 487248
rect 345018 487192 345074 487248
rect 349158 487192 349214 487248
rect 354678 487192 354734 487248
rect 360198 487192 360254 487248
rect 407946 636384 408002 636440
rect 407670 635296 407726 635352
rect 407578 627952 407634 628008
rect 407762 629584 407818 629640
rect 407670 526496 407726 526552
rect 407670 523232 407726 523288
rect 407578 520920 407634 520976
rect 407394 517928 407450 517984
rect 407854 607688 407910 607744
rect 407762 520240 407818 520296
rect 408130 633664 408186 633720
rect 408038 632576 408094 632632
rect 407854 498344 407910 498400
rect 408222 630944 408278 631000
rect 408314 610000 408370 610056
rect 408038 523232 408094 523288
rect 408038 498208 408094 498264
rect 407578 488280 407634 488336
rect 407394 488144 407450 488200
rect 408406 608640 408462 608696
rect 408314 500248 408370 500304
rect 408406 498616 408462 498672
rect 408406 498208 408462 498264
rect 440238 597488 440294 597544
rect 449898 597488 449954 597544
rect 459558 597488 459614 597544
rect 427818 597352 427874 597408
rect 430578 597352 430634 597408
rect 434718 597352 434774 597408
rect 422574 597216 422630 597272
rect 426438 597216 426494 597272
rect 409326 596808 409382 596864
rect 423678 596944 423734 597000
rect 429198 596944 429254 597000
rect 433338 597080 433394 597136
rect 434718 597100 434774 597136
rect 434718 597080 434720 597100
rect 434720 597080 434772 597100
rect 434772 597080 434774 597100
rect 431958 596944 432014 597000
rect 434718 596672 434774 596728
rect 425058 596420 425114 596456
rect 425058 596400 425060 596420
rect 425060 596400 425112 596420
rect 425112 596400 425114 596420
rect 444378 596672 444434 596728
rect 455418 596264 455474 596320
rect 470598 596264 470654 596320
rect 470598 589872 470654 589928
rect 422574 488416 422630 488472
rect 423678 488436 423734 488472
rect 423678 488416 423680 488436
rect 423680 488416 423732 488436
rect 423732 488416 423734 488436
rect 425058 488452 425060 488472
rect 425060 488452 425112 488472
rect 425112 488452 425114 488472
rect 425058 488416 425114 488452
rect 465078 488280 465134 488336
rect 429198 488144 429254 488200
rect 434718 488144 434774 488200
rect 426438 487600 426494 487656
rect 427818 487620 427874 487656
rect 427818 487600 427820 487620
rect 427820 487600 427872 487620
rect 427872 487600 427874 487620
rect 430578 487736 430634 487792
rect 433338 487464 433394 487520
rect 432142 487328 432198 487384
rect 434718 487348 434774 487384
rect 434718 487328 434720 487348
rect 434720 487328 434772 487348
rect 434772 487328 434774 487348
rect 434718 487192 434774 487248
rect 440238 487192 440294 487248
rect 444378 487192 444434 487248
rect 449898 487192 449954 487248
rect 455418 487192 455474 487248
rect 459558 487192 459614 487248
rect 470598 487192 470654 487248
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 299386 448568 299442 448624
rect 298834 446256 298890 446312
rect 296810 439456 296866 439512
rect 296902 434696 296958 434752
rect 298006 443536 298062 443592
rect 298006 430616 298062 430672
rect 298006 425856 298062 425912
rect 297638 421776 297694 421832
rect 297546 417016 297602 417072
rect 297454 412936 297510 412992
rect 297362 408176 297418 408232
rect 298006 404096 298062 404152
rect 298742 443808 298798 443864
rect 292578 6568 292634 6624
rect 298926 443128 298982 443184
rect 299110 443264 299166 443320
rect 299294 443400 299350 443456
rect 383934 454008 383990 454064
rect 384026 452240 384082 452296
rect 384026 448160 384082 448216
rect 383934 438640 383990 438696
rect 383934 421640 383990 421696
rect 385314 442856 385370 442912
rect 385222 434016 385278 434072
rect 580170 431568 580226 431624
rect 385130 429936 385186 429992
rect 580262 418240 580318 418296
rect 385038 416336 385094 416392
rect 385038 407496 385094 407552
rect 579986 404912 580042 404968
rect 382738 400696 382794 400752
rect 390558 400288 390614 400344
rect 316130 398520 316186 398576
rect 329010 399064 329066 399120
rect 337382 398792 337438 398848
rect 374734 398656 374790 398712
rect 379242 397840 379298 397896
rect 310518 397296 310574 397352
rect 307758 25472 307814 25528
rect 303158 3984 303214 4040
rect 307850 18536 307906 18592
rect 324318 397160 324374 397216
rect 310242 7656 310298 7712
rect 313830 3848 313886 3904
rect 364338 397024 364394 397080
rect 328458 83408 328514 83464
rect 326802 9016 326858 9072
rect 327998 7520 328054 7576
rect 343638 26968 343694 27024
rect 346398 19896 346454 19952
rect 339866 6296 339922 6352
rect 338670 3712 338726 3768
rect 345754 6432 345810 6488
rect 360198 352824 360254 352880
rect 361578 26832 361634 26888
rect 363510 8880 363566 8936
rect 378138 21664 378194 21720
rect 381174 10512 381230 10568
rect 382370 21528 382426 21584
rect 398838 396888 398894 396944
rect 398930 351056 398986 351112
rect 431958 396752 432014 396808
rect 414018 21392 414074 21448
rect 416778 21256 416834 21312
rect 412638 10376 412694 10432
rect 415398 10240 415454 10296
rect 434718 177248 434774 177304
rect 432050 16224 432106 16280
rect 433982 11736 434038 11792
rect 489918 398248 489974 398304
rect 452658 396616 452714 396672
rect 451646 11600 451702 11656
rect 470598 82048 470654 82104
rect 466458 22752 466514 22808
rect 469862 13096 469918 13152
rect 483018 397432 483074 397488
rect 488538 354184 488594 354240
rect 485778 22616 485834 22672
rect 484766 12960 484822 13016
rect 487618 3576 487674 3632
rect 494058 398112 494114 398168
rect 507858 397976 507914 398032
rect 506478 352688 506534 352744
rect 503718 24248 503774 24304
rect 505374 3440 505430 3496
rect 521658 395392 521714 395448
rect 520278 14456 520334 14512
rect 523774 16088 523830 16144
rect 523038 4936 523094 4992
rect 538218 354048 538274 354104
rect 539598 86128 539654 86184
rect 541990 15952 542046 16008
rect 540794 4800 540850 4856
rect 556158 395256 556214 395312
rect 557538 355272 557594 355328
rect 558918 353912 558974 353968
rect 556250 15816 556306 15872
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 576858 352552 576914 352608
rect 574098 24112 574154 24168
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 576306 6160 576362 6216
rect 579802 3304 579858 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3601 658202 3667 658205
rect -960 658200 3667 658202
rect -960 658144 3606 658200
rect 3662 658144 3667 658200
rect -960 658142 3667 658144
rect -960 658052 480 658142
rect 3601 658139 3667 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 187325 637122 187391 637125
rect 187325 637120 189458 637122
rect 187325 637064 187330 637120
rect 187386 637064 189458 637120
rect 187325 637062 189458 637064
rect 187325 637059 187391 637062
rect 189398 637060 189458 637062
rect 78581 636442 78647 636445
rect 80002 636442 80062 637030
rect 189398 637000 190072 637060
rect 299430 637000 300012 637060
rect 298001 636986 298067 636989
rect 299430 636986 299490 637000
rect 298001 636984 299490 636986
rect 298001 636928 298006 636984
rect 298062 636928 299490 636984
rect 298001 636926 299490 636928
rect 298001 636923 298067 636926
rect 78581 636440 80062 636442
rect 78581 636384 78586 636440
rect 78642 636384 80062 636440
rect 78581 636382 80062 636384
rect 407941 636442 408007 636445
rect 410002 636442 410062 637030
rect 407941 636440 410062 636442
rect 407941 636384 407946 636440
rect 408002 636384 410062 636440
rect 407941 636382 410062 636384
rect 78581 636379 78647 636382
rect 407941 636379 408007 636382
rect 186773 636034 186839 636037
rect 186773 636032 189458 636034
rect 186773 635976 186778 636032
rect 186834 635976 189458 636032
rect 186773 635974 189458 635976
rect 186773 635971 186839 635974
rect 189398 635972 189458 635974
rect 78305 635354 78371 635357
rect 80002 635354 80062 635942
rect 189398 635912 190072 635972
rect 299430 635912 300012 635972
rect 297173 635898 297239 635901
rect 299430 635898 299490 635912
rect 297173 635896 299490 635898
rect 297173 635840 297178 635896
rect 297234 635840 299490 635896
rect 297173 635838 299490 635840
rect 297173 635835 297239 635838
rect 78305 635352 80062 635354
rect 78305 635296 78310 635352
rect 78366 635296 80062 635352
rect 78305 635294 80062 635296
rect 407665 635354 407731 635357
rect 410002 635354 410062 635942
rect 407665 635352 410062 635354
rect 407665 635296 407670 635352
rect 407726 635296 410062 635352
rect 407665 635294 410062 635296
rect 78305 635291 78371 635294
rect 407665 635291 407731 635294
rect 186865 634402 186931 634405
rect 186865 634400 189458 634402
rect 186865 634344 186870 634400
rect 186926 634344 189458 634400
rect 186865 634342 189458 634344
rect 186865 634339 186931 634342
rect 189398 634340 189458 634342
rect 78213 633722 78279 633725
rect 80002 633722 80062 634310
rect 189398 634280 190072 634340
rect 299430 634280 300012 634340
rect 297909 634266 297975 634269
rect 299430 634266 299490 634280
rect 297909 634264 299490 634266
rect 297909 634208 297914 634264
rect 297970 634208 299490 634264
rect 297909 634206 299490 634208
rect 297909 634203 297975 634206
rect 78213 633720 80062 633722
rect 78213 633664 78218 633720
rect 78274 633664 80062 633720
rect 78213 633662 80062 633664
rect 408125 633722 408191 633725
rect 410002 633722 410062 634310
rect 408125 633720 410062 633722
rect 408125 633664 408130 633720
rect 408186 633664 410062 633720
rect 408125 633662 410062 633664
rect 78213 633659 78279 633662
rect 408125 633659 408191 633662
rect 187417 633314 187483 633317
rect 187417 633312 189458 633314
rect 187417 633256 187422 633312
rect 187478 633256 189458 633312
rect 187417 633254 189458 633256
rect 187417 633251 187483 633254
rect 189398 633252 189458 633254
rect 77753 632634 77819 632637
rect 80002 632634 80062 633222
rect 189398 633192 190072 633252
rect 299430 633192 300012 633252
rect 297725 633178 297791 633181
rect 299430 633178 299490 633192
rect 297725 633176 299490 633178
rect 297725 633120 297730 633176
rect 297786 633120 299490 633176
rect 297725 633118 299490 633120
rect 297725 633115 297791 633118
rect 77753 632632 80062 632634
rect 77753 632576 77758 632632
rect 77814 632576 80062 632632
rect 77753 632574 80062 632576
rect 408033 632634 408099 632637
rect 410002 632634 410062 633222
rect 408033 632632 410062 632634
rect 408033 632576 408038 632632
rect 408094 632576 410062 632632
rect 408033 632574 410062 632576
rect 77753 632571 77819 632574
rect 408033 632571 408099 632574
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 187233 631682 187299 631685
rect 187233 631680 189458 631682
rect 187233 631624 187238 631680
rect 187294 631624 189458 631680
rect 187233 631622 189458 631624
rect 187233 631619 187299 631622
rect 189398 631620 189458 631622
rect 78121 631002 78187 631005
rect 80002 631002 80062 631590
rect 189398 631560 190072 631620
rect 299430 631560 300012 631620
rect 297449 631546 297515 631549
rect 299430 631546 299490 631560
rect 297449 631544 299490 631546
rect 297449 631488 297454 631544
rect 297510 631488 299490 631544
rect 297449 631486 299490 631488
rect 297449 631483 297515 631486
rect 78121 631000 80062 631002
rect 78121 630944 78126 631000
rect 78182 630944 80062 631000
rect 78121 630942 80062 630944
rect 408217 631002 408283 631005
rect 410002 631002 410062 631590
rect 408217 631000 410062 631002
rect 408217 630944 408222 631000
rect 408278 630944 410062 631000
rect 408217 630942 410062 630944
rect 78121 630939 78187 630942
rect 408217 630939 408283 630942
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect 187509 630322 187575 630325
rect 187509 630320 189458 630322
rect 187509 630264 187514 630320
rect 187570 630264 189458 630320
rect 187509 630262 189458 630264
rect 187509 630259 187575 630262
rect 189398 630260 189458 630262
rect 77845 629642 77911 629645
rect 80002 629642 80062 630230
rect 189398 630200 190072 630260
rect 299430 630200 300012 630260
rect 297817 630186 297883 630189
rect 299430 630186 299490 630200
rect 297817 630184 299490 630186
rect 297817 630128 297822 630184
rect 297878 630128 299490 630184
rect 297817 630126 299490 630128
rect 297817 630123 297883 630126
rect 77845 629640 80062 629642
rect 77845 629584 77850 629640
rect 77906 629584 80062 629640
rect 77845 629582 80062 629584
rect 407757 629642 407823 629645
rect 410002 629642 410062 630230
rect 407757 629640 410062 629642
rect 407757 629584 407762 629640
rect 407818 629584 410062 629640
rect 407757 629582 410062 629584
rect 77845 629579 77911 629582
rect 407757 629579 407823 629582
rect 187141 628690 187207 628693
rect 187141 628688 189458 628690
rect 187141 628632 187146 628688
rect 187202 628632 189458 628688
rect 187141 628630 189458 628632
rect 187141 628627 187207 628630
rect 189398 628628 189458 628630
rect 78029 628010 78095 628013
rect 80002 628010 80062 628598
rect 189398 628568 190072 628628
rect 299430 628568 300012 628628
rect 297541 628554 297607 628557
rect 299430 628554 299490 628568
rect 297541 628552 299490 628554
rect 297541 628496 297546 628552
rect 297602 628496 299490 628552
rect 297541 628494 299490 628496
rect 297541 628491 297607 628494
rect 78029 628008 80062 628010
rect 78029 627952 78034 628008
rect 78090 627952 80062 628008
rect 78029 627950 80062 627952
rect 407573 628010 407639 628013
rect 410002 628010 410062 628598
rect 407573 628008 410062 628010
rect 407573 627952 407578 628008
rect 407634 627952 410062 628008
rect 407573 627950 410062 627952
rect 78029 627947 78095 627950
rect 407573 627947 407639 627950
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 187049 610330 187115 610333
rect 187049 610328 189458 610330
rect 187049 610272 187054 610328
rect 187110 610272 189458 610328
rect 187049 610270 189458 610272
rect 187049 610267 187115 610270
rect 189398 610268 189458 610270
rect 78397 610058 78463 610061
rect 80002 610058 80062 610238
rect 189398 610208 190072 610268
rect 299430 610208 300012 610268
rect 297081 610194 297147 610197
rect 299430 610194 299490 610208
rect 297081 610192 299490 610194
rect 297081 610136 297086 610192
rect 297142 610136 299490 610192
rect 297081 610134 299490 610136
rect 297081 610131 297147 610134
rect 78397 610056 80062 610058
rect 78397 610000 78402 610056
rect 78458 610000 80062 610056
rect 78397 609998 80062 610000
rect 408309 610058 408375 610061
rect 410002 610058 410062 610238
rect 408309 610056 410062 610058
rect 408309 610000 408314 610056
rect 408370 610000 410062 610056
rect 408309 609998 410062 610000
rect 78397 609995 78463 609998
rect 408309 609995 408375 609998
rect 77937 608698 78003 608701
rect 187601 608698 187667 608701
rect 296989 608698 297055 608701
rect 408401 608698 408467 608701
rect 77937 608696 80062 608698
rect 77937 608640 77942 608696
rect 77998 608640 80062 608696
rect 77937 608638 80062 608640
rect 77937 608635 78003 608638
rect 80002 608606 80062 608638
rect 187601 608696 189458 608698
rect 187601 608640 187606 608696
rect 187662 608640 189458 608696
rect 187601 608638 189458 608640
rect 187601 608635 187667 608638
rect 189398 608636 189458 608638
rect 296989 608696 299490 608698
rect 296989 608640 296994 608696
rect 297050 608640 299490 608696
rect 296989 608638 299490 608640
rect 189398 608576 190072 608636
rect 296989 608635 297055 608638
rect 299430 608636 299490 608638
rect 408401 608696 410062 608698
rect 408401 608640 408406 608696
rect 408462 608640 410062 608696
rect 408401 608638 410062 608640
rect 299430 608576 300012 608636
rect 408401 608635 408467 608638
rect 410002 608606 410062 608638
rect 186957 608426 187023 608429
rect 186957 608424 189458 608426
rect 186957 608368 186962 608424
rect 187018 608368 189458 608424
rect 186957 608366 189458 608368
rect 186957 608363 187023 608366
rect 189398 608364 189458 608366
rect 78489 607746 78555 607749
rect 80002 607746 80062 608334
rect 189398 608304 190072 608364
rect 299430 608304 300012 608364
rect 297633 608290 297699 608293
rect 299430 608290 299490 608304
rect 297633 608288 299490 608290
rect 297633 608232 297638 608288
rect 297694 608232 299490 608288
rect 297633 608230 299490 608232
rect 297633 608227 297699 608230
rect 78489 607744 80062 607746
rect 78489 607688 78494 607744
rect 78550 607688 80062 607744
rect 78489 607686 80062 607688
rect 407849 607746 407915 607749
rect 410002 607746 410062 608334
rect 407849 607744 410062 607746
rect 407849 607688 407854 607744
rect 407910 607688 410062 607744
rect 407849 607686 410062 607688
rect 78489 607683 78555 607686
rect 407849 607683 407915 607686
rect -960 606114 480 606204
rect 3877 606114 3943 606117
rect -960 606112 3943 606114
rect -960 606056 3882 606112
rect 3938 606056 3943 606112
rect -960 606054 3943 606056
rect -960 605964 480 606054
rect 3877 606051 3943 606054
rect 583520 604060 584960 604300
rect 102358 597484 102364 597548
rect 102428 597546 102434 597548
rect 102869 597546 102935 597549
rect 102428 597544 102935 597546
rect 102428 597488 102874 597544
rect 102930 597488 102935 597544
rect 102428 597486 102935 597488
rect 102428 597484 102434 597486
rect 102869 597483 102935 597486
rect 110454 597484 110460 597548
rect 110524 597546 110530 597548
rect 111701 597546 111767 597549
rect 207841 597548 207907 597549
rect 208945 597548 209011 597549
rect 207790 597546 207796 597548
rect 110524 597544 111767 597546
rect 110524 597488 111706 597544
rect 111762 597488 111767 597544
rect 110524 597486 111767 597488
rect 207750 597486 207796 597546
rect 207860 597544 207907 597548
rect 208894 597546 208900 597548
rect 207902 597488 207907 597544
rect 110524 597484 110530 597486
rect 111701 597483 111767 597486
rect 207790 597484 207796 597486
rect 207860 597484 207907 597488
rect 208854 597486 208900 597546
rect 208964 597544 209011 597548
rect 209006 597488 209011 597544
rect 208894 597484 208900 597486
rect 208964 597484 209011 597488
rect 207841 597483 207907 597484
rect 208945 597483 209011 597484
rect 209957 597548 210023 597549
rect 211153 597548 211219 597549
rect 209957 597544 210004 597548
rect 210068 597546 210074 597548
rect 211102 597546 211108 597548
rect 209957 597488 209962 597544
rect 209957 597484 210004 597488
rect 210068 597486 210114 597546
rect 211062 597486 211108 597546
rect 211172 597544 211219 597548
rect 211214 597488 211219 597544
rect 210068 597484 210074 597486
rect 211102 597484 211108 597486
rect 211172 597484 211219 597488
rect 209957 597483 210023 597484
rect 211153 597483 211219 597484
rect 212349 597548 212415 597549
rect 212349 597544 212396 597548
rect 212460 597546 212466 597548
rect 212349 597488 212354 597544
rect 212349 597484 212396 597488
rect 212460 597486 212506 597546
rect 212460 597484 212466 597486
rect 213494 597484 213500 597548
rect 213564 597546 213570 597548
rect 213821 597546 213887 597549
rect 214833 597548 214899 597549
rect 214782 597546 214788 597548
rect 213564 597544 213887 597546
rect 213564 597488 213826 597544
rect 213882 597488 213887 597544
rect 213564 597486 213887 597488
rect 214742 597486 214788 597546
rect 214852 597544 214899 597548
rect 215293 597548 215359 597549
rect 215753 597548 215819 597549
rect 215293 597546 215340 597548
rect 214894 597488 214899 597544
rect 213564 597484 213570 597486
rect 212349 597483 212415 597484
rect 213821 597483 213887 597486
rect 214782 597484 214788 597486
rect 214852 597484 214899 597488
rect 215248 597544 215340 597546
rect 215248 597488 215298 597544
rect 215248 597486 215340 597488
rect 214833 597483 214899 597484
rect 215293 597484 215340 597486
rect 215404 597484 215410 597548
rect 215702 597546 215708 597548
rect 215662 597486 215708 597546
rect 215772 597544 215819 597548
rect 215814 597488 215819 597544
rect 215702 597484 215708 597486
rect 215772 597484 215819 597488
rect 225454 597484 225460 597548
rect 225524 597546 225530 597548
rect 226241 597546 226307 597549
rect 225524 597544 226307 597546
rect 225524 597488 226246 597544
rect 226302 597488 226307 597544
rect 225524 597486 226307 597488
rect 225524 597484 225530 597486
rect 215293 597483 215359 597484
rect 215753 597483 215819 597484
rect 226241 597483 226307 597486
rect 235574 597484 235580 597548
rect 235644 597546 235650 597548
rect 235901 597546 235967 597549
rect 245561 597548 245627 597549
rect 235644 597544 235967 597546
rect 235644 597488 235906 597544
rect 235962 597488 235967 597544
rect 235644 597486 235967 597488
rect 235644 597484 235650 597486
rect 235901 597483 235967 597486
rect 245510 597484 245516 597548
rect 245580 597546 245627 597548
rect 245580 597544 245672 597546
rect 245622 597488 245672 597544
rect 245580 597486 245672 597488
rect 245580 597484 245627 597486
rect 250478 597484 250484 597548
rect 250548 597546 250554 597548
rect 251081 597546 251147 597549
rect 317689 597548 317755 597549
rect 320081 597548 320147 597549
rect 317638 597546 317644 597548
rect 250548 597544 251147 597546
rect 250548 597488 251086 597544
rect 251142 597488 251147 597544
rect 250548 597486 251147 597488
rect 317598 597486 317644 597546
rect 317708 597544 317755 597548
rect 320030 597546 320036 597548
rect 317750 597488 317755 597544
rect 250548 597484 250554 597486
rect 245561 597483 245627 597484
rect 251081 597483 251147 597486
rect 317638 597484 317644 597486
rect 317708 597484 317755 597488
rect 319990 597486 320036 597546
rect 320100 597544 320147 597548
rect 320142 597488 320147 597544
rect 320030 597484 320036 597486
rect 320100 597484 320147 597488
rect 317689 597483 317755 597484
rect 320081 597483 320147 597484
rect 320909 597546 320975 597549
rect 322197 597548 322263 597549
rect 321134 597546 321140 597548
rect 320909 597544 321140 597546
rect 320909 597488 320914 597544
rect 320970 597488 321140 597544
rect 320909 597486 321140 597488
rect 320909 597483 320975 597486
rect 321134 597484 321140 597486
rect 321204 597484 321210 597548
rect 322197 597544 322244 597548
rect 322308 597546 322314 597548
rect 322933 597546 322999 597549
rect 323342 597546 323348 597548
rect 322197 597488 322202 597544
rect 322197 597484 322244 597488
rect 322308 597486 322354 597546
rect 322933 597544 323348 597546
rect 322933 597488 322938 597544
rect 322994 597488 323348 597544
rect 322933 597486 323348 597488
rect 322308 597484 322314 597486
rect 322197 597483 322263 597484
rect 322933 597483 322999 597486
rect 323342 597484 323348 597486
rect 323412 597484 323418 597548
rect 324313 597546 324379 597549
rect 325182 597546 325188 597548
rect 324313 597544 325188 597546
rect 324313 597488 324318 597544
rect 324374 597488 325188 597544
rect 324313 597486 325188 597488
rect 324313 597483 324379 597486
rect 325182 597484 325188 597486
rect 325252 597484 325258 597548
rect 325734 597484 325740 597548
rect 325804 597546 325810 597548
rect 326153 597546 326219 597549
rect 325804 597544 326219 597546
rect 325804 597488 326158 597544
rect 326214 597488 326219 597544
rect 325804 597486 326219 597488
rect 325804 597484 325810 597486
rect 326153 597483 326219 597486
rect 329833 597546 329899 597549
rect 330518 597546 330524 597548
rect 329833 597544 330524 597546
rect 329833 597488 329838 597544
rect 329894 597488 330524 597544
rect 329833 597486 330524 597488
rect 329833 597483 329899 597486
rect 330518 597484 330524 597486
rect 330588 597484 330594 597548
rect 345013 597546 345079 597549
rect 345606 597546 345612 597548
rect 345013 597544 345612 597546
rect 345013 597488 345018 597544
rect 345074 597488 345612 597544
rect 345013 597486 345612 597488
rect 345013 597483 345079 597486
rect 345606 597484 345612 597486
rect 345676 597484 345682 597548
rect 360193 597546 360259 597549
rect 360510 597546 360516 597548
rect 360193 597544 360516 597546
rect 360193 597488 360198 597544
rect 360254 597488 360516 597544
rect 360193 597486 360516 597488
rect 360193 597483 360259 597486
rect 360510 597484 360516 597486
rect 360580 597484 360586 597548
rect 440233 597546 440299 597549
rect 440366 597546 440372 597548
rect 440233 597544 440372 597546
rect 440233 597488 440238 597544
rect 440294 597488 440372 597544
rect 440233 597486 440372 597488
rect 440233 597483 440299 597486
rect 440366 597484 440372 597486
rect 440436 597484 440442 597548
rect 449893 597546 449959 597549
rect 450486 597546 450492 597548
rect 449893 597544 450492 597546
rect 449893 597488 449898 597544
rect 449954 597488 450492 597544
rect 449893 597486 450492 597488
rect 449893 597483 449959 597486
rect 450486 597484 450492 597486
rect 450556 597484 450562 597548
rect 459553 597546 459619 597549
rect 460422 597546 460428 597548
rect 459553 597544 460428 597546
rect 459553 597488 459558 597544
rect 459614 597488 460428 597544
rect 459553 597486 460428 597488
rect 459553 597483 459619 597486
rect 460422 597484 460428 597486
rect 460492 597484 460498 597548
rect 92473 597410 92539 597413
rect 92974 597410 92980 597412
rect 92473 597408 92980 597410
rect 92473 597352 92478 597408
rect 92534 597352 92980 597408
rect 92473 597350 92980 597352
rect 92473 597347 92539 597350
rect 92974 597348 92980 597350
rect 93044 597348 93050 597412
rect 99966 597348 99972 597412
rect 100036 597410 100042 597412
rect 100661 597410 100727 597413
rect 100036 597408 100727 597410
rect 100036 597352 100666 597408
rect 100722 597352 100727 597408
rect 100036 597350 100727 597352
rect 100036 597348 100042 597350
rect 100661 597347 100727 597350
rect 318926 597348 318932 597412
rect 318996 597410 319002 597412
rect 319989 597410 320055 597413
rect 318996 597408 320055 597410
rect 318996 597352 319994 597408
rect 320050 597352 320055 597408
rect 318996 597350 320055 597352
rect 318996 597348 319002 597350
rect 319989 597347 320055 597350
rect 324405 597410 324471 597413
rect 324814 597410 324820 597412
rect 324405 597408 324820 597410
rect 324405 597352 324410 597408
rect 324466 597352 324820 597408
rect 324405 597350 324820 597352
rect 324405 597347 324471 597350
rect 324814 597348 324820 597350
rect 324884 597348 324890 597412
rect 335118 597348 335124 597412
rect 335188 597410 335194 597412
rect 335353 597410 335419 597413
rect 335188 597408 335419 597410
rect 335188 597352 335358 597408
rect 335414 597352 335419 597408
rect 335188 597350 335419 597352
rect 335188 597348 335194 597350
rect 335353 597347 335419 597350
rect 427813 597410 427879 597413
rect 428958 597410 428964 597412
rect 427813 597408 428964 597410
rect 427813 597352 427818 597408
rect 427874 597352 428964 597408
rect 427813 597350 428964 597352
rect 427813 597347 427879 597350
rect 428958 597348 428964 597350
rect 429028 597348 429034 597412
rect 430573 597410 430639 597413
rect 430982 597410 430988 597412
rect 430573 597408 430988 597410
rect 430573 597352 430578 597408
rect 430634 597352 430988 597408
rect 430573 597350 430988 597352
rect 430573 597347 430639 597350
rect 430982 597348 430988 597350
rect 431052 597348 431058 597412
rect 434713 597410 434779 597413
rect 435582 597410 435588 597412
rect 434713 597408 435588 597410
rect 434713 597352 434718 597408
rect 434774 597352 435588 597408
rect 434713 597350 435588 597352
rect 434713 597347 434779 597350
rect 435582 597348 435588 597350
rect 435652 597348 435658 597412
rect 98862 597212 98868 597276
rect 98932 597274 98938 597276
rect 99281 597274 99347 597277
rect 104801 597276 104867 597277
rect 98932 597272 99347 597274
rect 98932 597216 99286 597272
rect 99342 597216 99347 597272
rect 98932 597214 99347 597216
rect 98932 597212 98938 597214
rect 99281 597211 99347 597214
rect 104750 597212 104756 597276
rect 104820 597274 104867 597276
rect 104820 597272 104912 597274
rect 104862 597216 104912 597272
rect 104820 597214 104912 597216
rect 104820 597212 104867 597214
rect 230606 597212 230612 597276
rect 230676 597274 230682 597276
rect 231761 597274 231827 597277
rect 230676 597272 231827 597274
rect 230676 597216 231766 597272
rect 231822 597216 231827 597272
rect 230676 597214 231827 597216
rect 230676 597212 230682 597214
rect 104801 597211 104867 597212
rect 231761 597211 231827 597214
rect 313273 597274 313339 597277
rect 314326 597274 314332 597276
rect 313273 597272 314332 597274
rect 313273 597216 313278 597272
rect 313334 597216 314332 597272
rect 313273 597214 314332 597216
rect 313273 597211 313339 597214
rect 314326 597212 314332 597214
rect 314396 597212 314402 597276
rect 422569 597274 422635 597277
rect 422886 597274 422892 597276
rect 422569 597272 422892 597274
rect 422569 597216 422574 597272
rect 422630 597216 422892 597272
rect 422569 597214 422892 597216
rect 422569 597211 422635 597214
rect 422886 597212 422892 597214
rect 422956 597212 422962 597276
rect 426433 597274 426499 597277
rect 427670 597274 427676 597276
rect 426433 597272 427676 597274
rect 426433 597216 426438 597272
rect 426494 597216 427676 597272
rect 426433 597214 427676 597216
rect 426433 597211 426499 597214
rect 427670 597212 427676 597214
rect 427740 597212 427746 597276
rect 94037 597138 94103 597141
rect 94262 597138 94268 597140
rect 94037 597136 94268 597138
rect 94037 597080 94042 597136
rect 94098 597080 94268 597136
rect 94037 597078 94268 597080
rect 94037 597075 94103 597078
rect 94262 597076 94268 597078
rect 94332 597076 94338 597140
rect 101070 597076 101076 597140
rect 101140 597138 101146 597140
rect 102041 597138 102107 597141
rect 101140 597136 102107 597138
rect 101140 597080 102046 597136
rect 102102 597080 102107 597136
rect 101140 597078 102107 597080
rect 101140 597076 101146 597078
rect 102041 597075 102107 597078
rect 204345 597138 204411 597141
rect 205398 597138 205404 597140
rect 204345 597136 205404 597138
rect 204345 597080 204350 597136
rect 204406 597080 205404 597136
rect 204345 597078 205404 597080
rect 204345 597075 204411 597078
rect 205398 597076 205404 597078
rect 205468 597076 205474 597140
rect 349153 597138 349219 597141
rect 433333 597140 433399 597141
rect 434713 597140 434779 597141
rect 350390 597138 350396 597140
rect 349153 597136 350396 597138
rect 349153 597080 349158 597136
rect 349214 597080 350396 597136
rect 349153 597078 350396 597080
rect 349153 597075 349219 597078
rect 350390 597076 350396 597078
rect 350460 597076 350466 597140
rect 433333 597138 433380 597140
rect 433288 597136 433380 597138
rect 433288 597080 433338 597136
rect 433288 597078 433380 597080
rect 433333 597076 433380 597078
rect 433444 597076 433450 597140
rect 434662 597076 434668 597140
rect 434732 597138 434779 597140
rect 434732 597136 434824 597138
rect 434774 597080 434824 597136
rect 434732 597078 434824 597080
rect 434732 597076 434779 597078
rect 433333 597075 433399 597076
rect 434713 597075 434779 597076
rect 103278 596940 103284 597004
rect 103348 597002 103354 597004
rect 103421 597002 103487 597005
rect 103348 597000 103487 597002
rect 103348 596944 103426 597000
rect 103482 596944 103487 597000
rect 103348 596942 103487 596944
rect 103348 596940 103354 596942
rect 103421 596939 103487 596942
rect 105670 596940 105676 597004
rect 105740 597002 105746 597004
rect 106181 597002 106247 597005
rect 105740 597000 106247 597002
rect 105740 596944 106186 597000
rect 106242 596944 106247 597000
rect 105740 596942 106247 596944
rect 105740 596940 105746 596942
rect 106181 596939 106247 596942
rect 130510 596940 130516 597004
rect 130580 597002 130586 597004
rect 131021 597002 131087 597005
rect 130580 597000 131087 597002
rect 130580 596944 131026 597000
rect 131082 596944 131087 597000
rect 130580 596942 131087 596944
rect 130580 596940 130586 596942
rect 131021 596939 131087 596942
rect 339493 597002 339559 597005
rect 340454 597002 340460 597004
rect 339493 597000 340460 597002
rect 339493 596944 339498 597000
rect 339554 596944 340460 597000
rect 339493 596942 340460 596944
rect 339493 596939 339559 596942
rect 340454 596940 340460 596942
rect 340524 596940 340530 597004
rect 423673 597002 423739 597005
rect 424174 597002 424180 597004
rect 423673 597000 424180 597002
rect 423673 596944 423678 597000
rect 423734 596944 424180 597000
rect 423673 596942 424180 596944
rect 423673 596939 423739 596942
rect 424174 596940 424180 596942
rect 424244 596940 424250 597004
rect 429193 597002 429259 597005
rect 429878 597002 429884 597004
rect 429193 597000 429884 597002
rect 429193 596944 429198 597000
rect 429254 596944 429884 597000
rect 429193 596942 429884 596944
rect 429193 596939 429259 596942
rect 429878 596940 429884 596942
rect 429948 596940 429954 597004
rect 431718 596940 431724 597004
rect 431788 597002 431794 597004
rect 431953 597002 432019 597005
rect 431788 597000 432019 597002
rect 431788 596944 431958 597000
rect 432014 596944 432019 597000
rect 431788 596942 432019 596944
rect 431788 596940 431794 596942
rect 431953 596939 432019 596942
rect 97758 596804 97764 596868
rect 97828 596866 97834 596868
rect 97901 596866 97967 596869
rect 97828 596864 97967 596866
rect 97828 596808 97906 596864
rect 97962 596808 97967 596864
rect 97828 596806 97967 596808
rect 97828 596804 97834 596806
rect 97901 596803 97967 596806
rect 105302 596804 105308 596868
rect 105372 596866 105378 596868
rect 173157 596866 173223 596869
rect 105372 596864 173223 596866
rect 105372 596808 173162 596864
rect 173218 596808 173223 596864
rect 105372 596806 173223 596808
rect 105372 596804 105378 596806
rect 173157 596803 173223 596806
rect 240542 596804 240548 596868
rect 240612 596866 240618 596868
rect 241421 596866 241487 596869
rect 240612 596864 241487 596866
rect 240612 596808 241426 596864
rect 241482 596808 241487 596864
rect 240612 596806 241487 596808
rect 240612 596804 240618 596806
rect 241421 596803 241487 596806
rect 314653 596866 314719 596869
rect 315246 596866 315252 596868
rect 314653 596864 315252 596866
rect 314653 596808 314658 596864
rect 314714 596808 315252 596864
rect 314653 596806 315252 596808
rect 314653 596803 314719 596806
rect 315246 596804 315252 596806
rect 315316 596804 315322 596868
rect 409321 596866 409387 596869
rect 465390 596866 465396 596868
rect 409321 596864 465396 596866
rect 409321 596808 409326 596864
rect 409382 596808 465396 596864
rect 409321 596806 465396 596808
rect 409321 596803 409387 596806
rect 465390 596804 465396 596806
rect 465460 596804 465466 596868
rect 125542 596668 125548 596732
rect 125612 596730 125618 596732
rect 126881 596730 126947 596733
rect 125612 596728 126947 596730
rect 125612 596672 126886 596728
rect 126942 596672 126947 596728
rect 125612 596670 126947 596672
rect 125612 596668 125618 596670
rect 126881 596667 126947 596670
rect 434713 596730 434779 596733
rect 435214 596730 435220 596732
rect 434713 596728 435220 596730
rect 434713 596672 434718 596728
rect 434774 596672 435220 596728
rect 434713 596670 435220 596672
rect 434713 596667 434779 596670
rect 435214 596668 435220 596670
rect 435284 596668 435290 596732
rect 444373 596730 444439 596733
rect 445518 596730 445524 596732
rect 444373 596728 445524 596730
rect 444373 596672 444378 596728
rect 444434 596672 445524 596728
rect 444373 596670 445524 596672
rect 444373 596667 444439 596670
rect 445518 596668 445524 596670
rect 445588 596668 445594 596732
rect 135478 596532 135484 596596
rect 135548 596594 135554 596596
rect 136541 596594 136607 596597
rect 140681 596596 140747 596597
rect 135548 596592 136607 596594
rect 135548 596536 136546 596592
rect 136602 596536 136607 596592
rect 135548 596534 136607 596536
rect 135548 596532 135554 596534
rect 136541 596531 136607 596534
rect 140630 596532 140636 596596
rect 140700 596594 140747 596596
rect 311893 596594 311959 596597
rect 312854 596594 312860 596596
rect 140700 596592 140792 596594
rect 140742 596536 140792 596592
rect 140700 596534 140792 596536
rect 311893 596592 312860 596594
rect 311893 596536 311898 596592
rect 311954 596536 312860 596592
rect 311893 596534 312860 596536
rect 140700 596532 140747 596534
rect 140681 596531 140747 596532
rect 311893 596531 311959 596534
rect 312854 596532 312860 596534
rect 312924 596532 312930 596596
rect 202873 596460 202939 596461
rect 202822 596396 202828 596460
rect 202892 596458 202939 596460
rect 425053 596458 425119 596461
rect 425278 596458 425284 596460
rect 202892 596456 202984 596458
rect 202934 596400 202984 596456
rect 202892 596398 202984 596400
rect 425053 596456 425284 596458
rect 425053 596400 425058 596456
rect 425114 596400 425284 596456
rect 425053 596398 425284 596400
rect 202892 596396 202939 596398
rect 202873 596395 202939 596396
rect 425053 596395 425119 596398
rect 425278 596396 425284 596398
rect 425348 596396 425354 596460
rect 95233 596322 95299 596325
rect 95366 596322 95372 596324
rect 95233 596320 95372 596322
rect 95233 596264 95238 596320
rect 95294 596264 95372 596320
rect 95233 596262 95372 596264
rect 95233 596259 95299 596262
rect 95366 596260 95372 596262
rect 95436 596260 95442 596324
rect 115606 596260 115612 596324
rect 115676 596322 115682 596324
rect 115841 596322 115907 596325
rect 115676 596320 115907 596322
rect 115676 596264 115846 596320
rect 115902 596264 115907 596320
rect 115676 596262 115907 596264
rect 115676 596260 115682 596262
rect 115841 596259 115907 596262
rect 120574 596260 120580 596324
rect 120644 596322 120650 596324
rect 121361 596322 121427 596325
rect 204253 596324 204319 596325
rect 204253 596322 204300 596324
rect 120644 596320 121427 596322
rect 120644 596264 121366 596320
rect 121422 596264 121427 596320
rect 120644 596262 121427 596264
rect 204208 596320 204300 596322
rect 204208 596264 204258 596320
rect 204208 596262 204300 596264
rect 120644 596260 120650 596262
rect 121361 596259 121427 596262
rect 204253 596260 204300 596262
rect 204364 596260 204370 596324
rect 219198 596260 219204 596324
rect 219268 596322 219274 596324
rect 219433 596322 219499 596325
rect 219268 596320 219499 596322
rect 219268 596264 219438 596320
rect 219494 596264 219499 596320
rect 219268 596262 219499 596264
rect 219268 596260 219274 596262
rect 204253 596259 204319 596260
rect 219433 596259 219499 596262
rect 354438 596260 354444 596324
rect 354508 596322 354514 596324
rect 354673 596322 354739 596325
rect 455413 596324 455479 596325
rect 455413 596322 455460 596324
rect 354508 596320 354739 596322
rect 354508 596264 354678 596320
rect 354734 596264 354739 596320
rect 354508 596262 354739 596264
rect 455368 596320 455460 596322
rect 455368 596264 455418 596320
rect 455368 596262 455460 596264
rect 354508 596260 354514 596262
rect 354673 596259 354739 596262
rect 455413 596260 455460 596262
rect 455524 596260 455530 596324
rect 470358 596260 470364 596324
rect 470428 596322 470434 596324
rect 470593 596322 470659 596325
rect 470428 596320 470659 596322
rect 470428 596264 470598 596320
rect 470654 596264 470659 596320
rect 470428 596262 470659 596264
rect 470428 596260 470434 596262
rect 455413 596259 455479 596260
rect 470593 596259 470659 596262
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 282126 589868 282132 589932
rect 282196 589930 282202 589932
rect 470593 589930 470659 589933
rect 282196 589928 470659 589930
rect 282196 589872 470598 589928
rect 470654 589872 470659 589928
rect 282196 589870 470659 589872
rect 282196 589868 282202 589870
rect 470593 589867 470659 589870
rect -960 580002 480 580092
rect 3969 580002 4035 580005
rect -960 580000 4035 580002
rect -960 579944 3974 580000
rect 4030 579944 4035 580000
rect -960 579942 4035 579944
rect -960 579852 480 579942
rect 3969 579939 4035 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 187325 527098 187391 527101
rect 298001 527098 298067 527101
rect 187325 527096 189458 527098
rect 187325 527040 187330 527096
rect 187386 527060 189458 527096
rect 298001 527096 299490 527098
rect 187386 527040 190072 527060
rect 187325 527038 190072 527040
rect 187325 527035 187391 527038
rect 78489 526690 78555 526693
rect 80002 526690 80062 527030
rect 189398 527000 190072 527038
rect 298001 527040 298006 527096
rect 298062 527060 299490 527096
rect 298062 527040 300012 527060
rect 298001 527038 300012 527040
rect 298001 527035 298067 527038
rect 299430 527000 300012 527038
rect 78489 526688 80062 526690
rect 78489 526632 78494 526688
rect 78550 526632 80062 526688
rect 78489 526630 80062 526632
rect 78489 526627 78555 526630
rect 407798 526628 407804 526692
rect 407868 526690 407874 526692
rect 410002 526690 410062 527030
rect 407868 526630 410062 526690
rect 407868 526628 407874 526630
rect 78305 526554 78371 526557
rect 407665 526554 407731 526557
rect 78305 526552 80062 526554
rect 78305 526496 78310 526552
rect 78366 526496 80062 526552
rect 78305 526494 80062 526496
rect 78305 526491 78371 526494
rect 80002 525942 80062 526494
rect 407665 526552 410062 526554
rect 407665 526496 407670 526552
rect 407726 526496 410062 526552
rect 407665 526494 410062 526496
rect 407665 526491 407731 526494
rect 186773 526010 186839 526013
rect 188429 526010 188495 526013
rect 297173 526010 297239 526013
rect 186773 526008 189458 526010
rect 186773 525952 186778 526008
rect 186834 525952 188434 526008
rect 188490 525972 189458 526008
rect 297173 526008 299490 526010
rect 188490 525952 190072 525972
rect 186773 525950 190072 525952
rect 186773 525947 186839 525950
rect 188429 525947 188495 525950
rect 189398 525912 190072 525950
rect 297173 525952 297178 526008
rect 297234 525972 299490 526008
rect 297234 525952 300012 525972
rect 297173 525950 300012 525952
rect 297173 525947 297239 525950
rect 299430 525912 300012 525950
rect 410002 525942 410062 526494
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 186865 524378 186931 524381
rect 187325 524378 187391 524381
rect 297357 524378 297423 524381
rect 297817 524378 297883 524381
rect 186865 524376 189458 524378
rect 186865 524320 186870 524376
rect 186926 524320 187330 524376
rect 187386 524340 189458 524376
rect 297357 524376 299490 524378
rect 187386 524320 190072 524340
rect 186865 524318 190072 524320
rect 186865 524315 186931 524318
rect 187325 524315 187391 524318
rect 78305 523698 78371 523701
rect 80002 523698 80062 524310
rect 189398 524280 190072 524318
rect 297357 524320 297362 524376
rect 297418 524320 297822 524376
rect 297878 524340 299490 524376
rect 583520 524364 584960 524454
rect 297878 524320 300012 524340
rect 297357 524318 300012 524320
rect 297357 524315 297423 524318
rect 297817 524315 297883 524318
rect 299430 524280 300012 524318
rect 78305 523696 80062 523698
rect 78305 523640 78310 523696
rect 78366 523640 80062 523696
rect 78305 523638 80062 523640
rect 78305 523635 78371 523638
rect 408166 523636 408172 523700
rect 408236 523698 408242 523700
rect 410002 523698 410062 524310
rect 408236 523638 410062 523698
rect 408236 523636 408242 523638
rect 77753 523562 77819 523565
rect 77753 523560 80062 523562
rect 77753 523504 77758 523560
rect 77814 523504 80062 523560
rect 77753 523502 80062 523504
rect 77753 523499 77819 523502
rect 80002 523222 80062 523502
rect 186773 523290 186839 523293
rect 187417 523290 187483 523293
rect 297725 523290 297791 523293
rect 407665 523290 407731 523293
rect 408033 523290 408099 523293
rect 186773 523288 189458 523290
rect 186773 523232 186778 523288
rect 186834 523232 187422 523288
rect 187478 523252 189458 523288
rect 297725 523288 299490 523290
rect 187478 523232 190072 523252
rect 186773 523230 190072 523232
rect 186773 523227 186839 523230
rect 187417 523227 187483 523230
rect 189398 523192 190072 523230
rect 297725 523232 297730 523288
rect 297786 523252 299490 523288
rect 407665 523288 410062 523290
rect 297786 523232 300012 523252
rect 297725 523230 300012 523232
rect 297725 523227 297791 523230
rect 299430 523192 300012 523230
rect 407665 523232 407670 523288
rect 407726 523232 408038 523288
rect 408094 523232 410062 523288
rect 407665 523230 410062 523232
rect 407665 523227 407731 523230
rect 408033 523227 408099 523230
rect 410002 523222 410062 523230
rect 77845 521658 77911 521661
rect 78121 521658 78187 521661
rect 77845 521656 78187 521658
rect 77845 521600 77850 521656
rect 77906 521600 78126 521656
rect 78182 521600 78187 521656
rect 77845 521598 78187 521600
rect 77845 521595 77911 521598
rect 78121 521595 78187 521598
rect 187233 521658 187299 521661
rect 297449 521658 297515 521661
rect 187233 521656 189458 521658
rect 187233 521600 187238 521656
rect 187294 521620 189458 521656
rect 297449 521656 299490 521658
rect 187294 521600 190072 521620
rect 187233 521598 190072 521600
rect 187233 521595 187299 521598
rect 77661 520978 77727 520981
rect 80002 520978 80062 521590
rect 189398 521560 190072 521598
rect 297449 521600 297454 521656
rect 297510 521620 299490 521656
rect 297510 521600 300012 521620
rect 297449 521598 300012 521600
rect 297449 521595 297515 521598
rect 299430 521560 300012 521598
rect 186865 521522 186931 521525
rect 187509 521522 187575 521525
rect 186865 521520 187575 521522
rect 186865 521464 186870 521520
rect 186926 521464 187514 521520
rect 187570 521464 187575 521520
rect 186865 521462 187575 521464
rect 186865 521459 186931 521462
rect 187509 521459 187575 521462
rect 77661 520976 80062 520978
rect 77661 520920 77666 520976
rect 77722 520920 80062 520976
rect 77661 520918 80062 520920
rect 407573 520978 407639 520981
rect 410002 520978 410062 521590
rect 407573 520976 410062 520978
rect 407573 520920 407578 520976
rect 407634 520920 410062 520976
rect 407573 520918 410062 520920
rect 77661 520915 77727 520918
rect 407573 520915 407639 520918
rect 78121 520298 78187 520301
rect 186865 520298 186931 520301
rect 298001 520298 298067 520301
rect 407757 520298 407823 520301
rect 78121 520296 80062 520298
rect 78121 520240 78126 520296
rect 78182 520240 80062 520296
rect 78121 520238 80062 520240
rect 78121 520235 78187 520238
rect 80002 520230 80062 520238
rect 186865 520296 190010 520298
rect 186865 520240 186870 520296
rect 186926 520260 190010 520296
rect 298001 520296 299858 520298
rect 186926 520240 190072 520260
rect 186865 520238 190072 520240
rect 186865 520235 186931 520238
rect 189950 520200 190072 520238
rect 298001 520240 298006 520296
rect 298062 520260 299858 520296
rect 407757 520296 410062 520298
rect 298062 520240 300012 520260
rect 298001 520238 300012 520240
rect 298001 520235 298067 520238
rect 299798 520200 300012 520238
rect 407757 520240 407762 520296
rect 407818 520240 410062 520296
rect 407757 520238 410062 520240
rect 407757 520235 407823 520238
rect 410002 520230 410062 520238
rect 187141 518666 187207 518669
rect 297541 518666 297607 518669
rect 187141 518664 189458 518666
rect 187141 518608 187146 518664
rect 187202 518628 189458 518664
rect 297541 518664 299490 518666
rect 187202 518608 190072 518628
rect 187141 518606 190072 518608
rect 187141 518603 187207 518606
rect 78581 517986 78647 517989
rect 80002 517986 80062 518598
rect 189398 518568 190072 518606
rect 297541 518608 297546 518664
rect 297602 518628 299490 518664
rect 297602 518608 300012 518628
rect 297541 518606 300012 518608
rect 297541 518603 297607 518606
rect 299430 518568 300012 518606
rect 78581 517984 80062 517986
rect 78581 517928 78586 517984
rect 78642 517928 80062 517984
rect 78581 517926 80062 517928
rect 407389 517986 407455 517989
rect 410002 517986 410062 518598
rect 407389 517984 410062 517986
rect 407389 517928 407394 517984
rect 407450 517928 410062 517984
rect 407389 517926 410062 517928
rect 78581 517923 78647 517926
rect 407389 517923 407455 517926
rect 296897 517578 296963 517581
rect 297541 517578 297607 517581
rect 296897 517576 297607 517578
rect 296897 517520 296902 517576
rect 296958 517520 297546 517576
rect 297602 517520 297607 517576
rect 296897 517518 297607 517520
rect 296897 517515 296963 517518
rect 297541 517515 297607 517518
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 187049 500306 187115 500309
rect 297081 500306 297147 500309
rect 408309 500306 408375 500309
rect 187049 500304 189458 500306
rect 187049 500248 187054 500304
rect 187110 500268 189458 500304
rect 297081 500304 299490 500306
rect 187110 500248 190072 500268
rect 187049 500246 190072 500248
rect 187049 500243 187115 500246
rect 78029 499898 78095 499901
rect 80002 499898 80062 500238
rect 189398 500208 190072 500246
rect 297081 500248 297086 500304
rect 297142 500268 299490 500304
rect 408309 500304 410062 500306
rect 297142 500248 300012 500268
rect 297081 500246 300012 500248
rect 297081 500243 297147 500246
rect 299430 500208 300012 500246
rect 408309 500248 408314 500304
rect 408370 500248 410062 500304
rect 408309 500246 410062 500248
rect 408309 500243 408375 500246
rect 410002 500238 410062 500246
rect 78029 499896 80062 499898
rect 78029 499840 78034 499896
rect 78090 499840 80062 499896
rect 78029 499838 80062 499840
rect 78029 499835 78095 499838
rect 77937 498674 78003 498677
rect 187601 498674 187667 498677
rect 189073 498674 189139 498677
rect 297817 498674 297883 498677
rect 408401 498674 408467 498677
rect 77937 498672 80062 498674
rect 77937 498616 77942 498672
rect 77998 498616 80062 498672
rect 77937 498614 80062 498616
rect 77937 498611 78003 498614
rect 80002 498606 80062 498614
rect 187601 498672 189458 498674
rect 187601 498616 187606 498672
rect 187662 498616 189078 498672
rect 189134 498636 189458 498672
rect 297817 498672 299490 498674
rect 189134 498616 190072 498636
rect 187601 498614 190072 498616
rect 187601 498611 187667 498614
rect 189073 498611 189139 498614
rect 189398 498576 190072 498614
rect 297817 498616 297822 498672
rect 297878 498636 299490 498672
rect 408401 498672 410062 498674
rect 297878 498616 300012 498636
rect 297817 498614 300012 498616
rect 297817 498611 297883 498614
rect 299430 498576 300012 498614
rect 408401 498616 408406 498672
rect 408462 498616 410062 498672
rect 408401 498614 410062 498616
rect 408401 498611 408467 498614
rect 410002 498606 410062 498614
rect 78397 498402 78463 498405
rect 297633 498402 297699 498405
rect 407849 498402 407915 498405
rect 78397 498400 79426 498402
rect 78397 498344 78402 498400
rect 78458 498364 79426 498400
rect 297633 498400 299490 498402
rect 78458 498344 80032 498364
rect 78397 498342 80032 498344
rect 78397 498339 78463 498342
rect 79366 498304 80032 498342
rect 189398 498304 190072 498364
rect 297633 498344 297638 498400
rect 297694 498364 299490 498400
rect 407849 498400 409522 498402
rect 297694 498344 300012 498364
rect 297633 498342 300012 498344
rect 297633 498339 297699 498342
rect 299430 498304 300012 498342
rect 407849 498344 407854 498400
rect 407910 498364 409522 498400
rect 407910 498344 410032 498364
rect 407849 498342 410032 498344
rect 407849 498339 407915 498342
rect 409462 498304 410032 498342
rect 186681 498266 186747 498269
rect 186957 498266 187023 498269
rect 189398 498266 189458 498304
rect 186681 498264 189458 498266
rect 186681 498208 186686 498264
rect 186742 498208 186962 498264
rect 187018 498208 189458 498264
rect 186681 498206 189458 498208
rect 408033 498266 408099 498269
rect 408401 498266 408467 498269
rect 408033 498264 408467 498266
rect 408033 498208 408038 498264
rect 408094 498208 408406 498264
rect 408462 498208 408467 498264
rect 408033 498206 408467 498208
rect 186681 498203 186747 498206
rect 186957 498203 187023 498206
rect 408033 498203 408099 498206
rect 408401 498203 408467 498206
rect 583520 497844 584960 498084
rect 297909 489834 297975 489837
rect 408166 489834 408172 489836
rect 297909 489832 408172 489834
rect 297909 489776 297914 489832
rect 297970 489776 408172 489832
rect 297909 489774 408172 489776
rect 297909 489771 297975 489774
rect 408166 489772 408172 489774
rect 408236 489772 408242 489836
rect -960 488596 480 488836
rect 92933 488476 92999 488477
rect 94221 488476 94287 488477
rect 95325 488476 95391 488477
rect 97809 488476 97875 488477
rect 98913 488476 98979 488477
rect 100017 488476 100083 488477
rect 101121 488476 101187 488477
rect 102409 488476 102475 488477
rect 104801 488476 104867 488477
rect 105721 488476 105787 488477
rect 92933 488472 92980 488476
rect 93044 488474 93050 488476
rect 92933 488416 92938 488472
rect 92933 488412 92980 488416
rect 93044 488414 93090 488474
rect 94221 488472 94268 488476
rect 94332 488474 94338 488476
rect 94221 488416 94226 488472
rect 93044 488412 93050 488414
rect 94221 488412 94268 488416
rect 94332 488414 94378 488474
rect 95325 488472 95372 488476
rect 95436 488474 95442 488476
rect 97758 488474 97764 488476
rect 95325 488416 95330 488472
rect 94332 488412 94338 488414
rect 95325 488412 95372 488416
rect 95436 488414 95482 488474
rect 97718 488414 97764 488474
rect 97828 488472 97875 488476
rect 98862 488474 98868 488476
rect 97870 488416 97875 488472
rect 95436 488412 95442 488414
rect 97758 488412 97764 488414
rect 97828 488412 97875 488416
rect 98822 488414 98868 488474
rect 98932 488472 98979 488476
rect 99966 488474 99972 488476
rect 98974 488416 98979 488472
rect 98862 488412 98868 488414
rect 98932 488412 98979 488416
rect 99926 488414 99972 488474
rect 100036 488472 100083 488476
rect 101070 488474 101076 488476
rect 100078 488416 100083 488472
rect 99966 488412 99972 488414
rect 100036 488412 100083 488416
rect 101030 488414 101076 488474
rect 101140 488472 101187 488476
rect 102358 488474 102364 488476
rect 101182 488416 101187 488472
rect 101070 488412 101076 488414
rect 101140 488412 101187 488416
rect 102318 488414 102364 488474
rect 102428 488472 102475 488476
rect 104750 488474 104756 488476
rect 102470 488416 102475 488472
rect 102358 488412 102364 488414
rect 102428 488412 102475 488416
rect 104710 488414 104756 488474
rect 104820 488472 104867 488476
rect 105670 488474 105676 488476
rect 104862 488416 104867 488472
rect 104750 488412 104756 488414
rect 104820 488412 104867 488416
rect 105630 488414 105676 488474
rect 105740 488472 105787 488476
rect 105782 488416 105787 488472
rect 105670 488412 105676 488414
rect 105740 488412 105787 488416
rect 204294 488412 204300 488476
rect 204364 488474 204370 488476
rect 204713 488474 204779 488477
rect 214833 488476 214899 488477
rect 214782 488474 214788 488476
rect 204364 488472 204779 488474
rect 204364 488416 204718 488472
rect 204774 488416 204779 488472
rect 204364 488414 204779 488416
rect 214742 488414 214788 488474
rect 214852 488472 214899 488476
rect 214894 488416 214899 488472
rect 204364 488412 204370 488414
rect 92933 488411 92999 488412
rect 94221 488411 94287 488412
rect 95325 488411 95391 488412
rect 97809 488411 97875 488412
rect 98913 488411 98979 488412
rect 100017 488411 100083 488412
rect 101121 488411 101187 488412
rect 102409 488411 102475 488412
rect 104801 488411 104867 488412
rect 105721 488411 105787 488412
rect 204713 488411 204779 488414
rect 214782 488412 214788 488414
rect 214852 488412 214899 488416
rect 214833 488411 214899 488412
rect 293309 488474 293375 488477
rect 293861 488474 293927 488477
rect 293309 488472 293927 488474
rect 293309 488416 293314 488472
rect 293370 488416 293866 488472
rect 293922 488416 293927 488472
rect 293309 488414 293927 488416
rect 293309 488411 293375 488414
rect 293861 488411 293927 488414
rect 297357 488474 297423 488477
rect 297817 488474 297883 488477
rect 314285 488476 314351 488477
rect 315389 488476 315455 488477
rect 297357 488472 302250 488474
rect 297357 488416 297362 488472
rect 297418 488416 297822 488472
rect 297878 488416 302250 488472
rect 297357 488414 302250 488416
rect 297357 488411 297423 488414
rect 297817 488411 297883 488414
rect 211153 488340 211219 488341
rect 211102 488338 211108 488340
rect 211062 488278 211108 488338
rect 211172 488336 211219 488340
rect 211214 488280 211219 488336
rect 211102 488276 211108 488278
rect 211172 488276 211219 488280
rect 213494 488276 213500 488340
rect 213564 488338 213570 488340
rect 213729 488338 213795 488341
rect 215753 488340 215819 488341
rect 215702 488338 215708 488340
rect 213564 488336 213795 488338
rect 213564 488280 213734 488336
rect 213790 488280 213795 488336
rect 213564 488278 213795 488280
rect 215662 488278 215708 488338
rect 215772 488336 215819 488340
rect 215814 488280 215819 488336
rect 213564 488276 213570 488278
rect 211153 488275 211219 488276
rect 213729 488275 213795 488278
rect 215702 488276 215708 488278
rect 215772 488276 215819 488280
rect 215753 488275 215819 488276
rect 296897 488338 296963 488341
rect 297357 488338 297423 488341
rect 302190 488338 302250 488414
rect 314285 488472 314332 488476
rect 314396 488474 314402 488476
rect 314285 488416 314290 488472
rect 314285 488412 314332 488416
rect 314396 488414 314442 488474
rect 315389 488472 315436 488476
rect 315500 488474 315506 488476
rect 422569 488474 422635 488477
rect 422886 488474 422892 488476
rect 315389 488416 315394 488472
rect 314396 488412 314402 488414
rect 315389 488412 315436 488416
rect 315500 488414 315546 488474
rect 422569 488472 422892 488474
rect 422569 488416 422574 488472
rect 422630 488416 422892 488472
rect 422569 488414 422892 488416
rect 315500 488412 315506 488414
rect 314285 488411 314351 488412
rect 315389 488411 315455 488412
rect 422569 488411 422635 488414
rect 422886 488412 422892 488414
rect 422956 488412 422962 488476
rect 423673 488474 423739 488477
rect 424174 488474 424180 488476
rect 423673 488472 424180 488474
rect 423673 488416 423678 488472
rect 423734 488416 424180 488472
rect 423673 488414 424180 488416
rect 423673 488411 423739 488414
rect 424174 488412 424180 488414
rect 424244 488412 424250 488476
rect 425053 488474 425119 488477
rect 425278 488474 425284 488476
rect 425053 488472 425284 488474
rect 425053 488416 425058 488472
rect 425114 488416 425284 488472
rect 425053 488414 425284 488416
rect 425053 488411 425119 488414
rect 425278 488412 425284 488414
rect 425348 488412 425354 488476
rect 407573 488338 407639 488341
rect 296897 488336 298938 488338
rect 296897 488280 296902 488336
rect 296958 488280 297362 488336
rect 297418 488280 298938 488336
rect 296897 488278 298938 488280
rect 302190 488336 407639 488338
rect 302190 488280 407578 488336
rect 407634 488280 407639 488336
rect 302190 488278 407639 488280
rect 296897 488275 296963 488278
rect 297357 488275 297423 488278
rect 105302 488140 105308 488204
rect 105372 488202 105378 488204
rect 105813 488202 105879 488205
rect 105372 488200 105879 488202
rect 105372 488144 105818 488200
rect 105874 488144 105879 488200
rect 105372 488142 105879 488144
rect 105372 488140 105378 488142
rect 105813 488139 105879 488142
rect 110454 488140 110460 488204
rect 110524 488202 110530 488204
rect 111701 488202 111767 488205
rect 110524 488200 111767 488202
rect 110524 488144 111706 488200
rect 111762 488144 111767 488200
rect 110524 488142 111767 488144
rect 110524 488140 110530 488142
rect 111701 488139 111767 488142
rect 202873 488202 202939 488205
rect 203006 488202 203012 488204
rect 202873 488200 203012 488202
rect 202873 488144 202878 488200
rect 202934 488144 203012 488200
rect 202873 488142 203012 488144
rect 202873 488139 202939 488142
rect 203006 488140 203012 488142
rect 203076 488140 203082 488204
rect 298878 488202 298938 488278
rect 407573 488275 407639 488278
rect 465073 488338 465139 488341
rect 465390 488338 465396 488340
rect 465073 488336 465396 488338
rect 465073 488280 465078 488336
rect 465134 488280 465396 488336
rect 465073 488278 465396 488280
rect 465073 488275 465139 488278
rect 465390 488276 465396 488278
rect 465460 488276 465466 488340
rect 407389 488202 407455 488205
rect 298878 488200 407455 488202
rect 298878 488144 407394 488200
rect 407450 488144 407455 488200
rect 298878 488142 407455 488144
rect 407389 488139 407455 488142
rect 429193 488202 429259 488205
rect 429878 488202 429884 488204
rect 429193 488200 429884 488202
rect 429193 488144 429198 488200
rect 429254 488144 429884 488200
rect 429193 488142 429884 488144
rect 429193 488139 429259 488142
rect 429878 488140 429884 488142
rect 429948 488140 429954 488204
rect 434713 488202 434779 488205
rect 435582 488202 435588 488204
rect 434713 488200 435588 488202
rect 434713 488144 434718 488200
rect 434774 488144 435588 488200
rect 434713 488142 435588 488144
rect 434713 488139 434779 488142
rect 435582 488140 435588 488142
rect 435652 488140 435658 488204
rect 293861 488066 293927 488069
rect 407798 488066 407804 488068
rect 293861 488064 407804 488066
rect 293861 488008 293866 488064
rect 293922 488008 407804 488064
rect 293861 488006 407804 488008
rect 293861 488003 293927 488006
rect 407798 488004 407804 488006
rect 407868 488004 407874 488068
rect 103278 487868 103284 487932
rect 103348 487930 103354 487932
rect 103421 487930 103487 487933
rect 103348 487928 103487 487930
rect 103348 487872 103426 487928
rect 103482 487872 103487 487928
rect 103348 487870 103487 487872
rect 103348 487868 103354 487870
rect 103421 487867 103487 487870
rect 208853 487932 208919 487933
rect 312997 487932 313063 487933
rect 208853 487928 208900 487932
rect 208964 487930 208970 487932
rect 208853 487872 208858 487928
rect 208853 487868 208900 487872
rect 208964 487870 209010 487930
rect 312997 487928 313044 487932
rect 313108 487930 313114 487932
rect 324405 487930 324471 487933
rect 324630 487930 324636 487932
rect 312997 487872 313002 487928
rect 208964 487868 208970 487870
rect 312997 487868 313044 487872
rect 313108 487870 313154 487930
rect 324405 487928 324636 487930
rect 324405 487872 324410 487928
rect 324466 487872 324636 487928
rect 324405 487870 324636 487872
rect 313108 487868 313114 487870
rect 208853 487867 208919 487868
rect 312997 487867 313063 487868
rect 324405 487867 324471 487870
rect 324630 487868 324636 487870
rect 324700 487868 324706 487932
rect 325734 487732 325740 487796
rect 325804 487794 325810 487796
rect 326613 487794 326679 487797
rect 325804 487792 326679 487794
rect 325804 487736 326618 487792
rect 326674 487736 326679 487792
rect 325804 487734 326679 487736
rect 325804 487732 325810 487734
rect 326613 487731 326679 487734
rect 430573 487794 430639 487797
rect 430982 487794 430988 487796
rect 430573 487792 430988 487794
rect 430573 487736 430578 487792
rect 430634 487736 430988 487792
rect 430573 487734 430988 487736
rect 430573 487731 430639 487734
rect 430982 487732 430988 487734
rect 431052 487732 431058 487796
rect 426433 487658 426499 487661
rect 427670 487658 427676 487660
rect 426433 487656 427676 487658
rect 426433 487600 426438 487656
rect 426494 487600 427676 487656
rect 426433 487598 427676 487600
rect 426433 487595 426499 487598
rect 427670 487596 427676 487598
rect 427740 487596 427746 487660
rect 427813 487658 427879 487661
rect 428958 487658 428964 487660
rect 427813 487656 428964 487658
rect 427813 487600 427818 487656
rect 427874 487600 428964 487656
rect 427813 487598 428964 487600
rect 427813 487595 427879 487598
rect 428958 487596 428964 487598
rect 429028 487596 429034 487660
rect 212206 487460 212212 487524
rect 212276 487522 212282 487524
rect 212349 487522 212415 487525
rect 212276 487520 212415 487522
rect 212276 487464 212354 487520
rect 212410 487464 212415 487520
rect 212276 487462 212415 487464
rect 212276 487460 212282 487462
rect 212349 487459 212415 487462
rect 319989 487524 320055 487525
rect 319989 487520 320036 487524
rect 320100 487522 320106 487524
rect 322933 487522 322999 487525
rect 433333 487524 433399 487525
rect 323342 487522 323348 487524
rect 319989 487464 319994 487520
rect 319989 487460 320036 487464
rect 320100 487462 320146 487522
rect 322933 487520 323348 487522
rect 322933 487464 322938 487520
rect 322994 487464 323348 487520
rect 322933 487462 323348 487464
rect 320100 487460 320106 487462
rect 319989 487459 320055 487460
rect 322933 487459 322999 487462
rect 323342 487460 323348 487462
rect 323412 487460 323418 487524
rect 433333 487522 433380 487524
rect 433288 487520 433380 487522
rect 433288 487464 433338 487520
rect 433288 487462 433380 487464
rect 433333 487460 433380 487462
rect 433444 487460 433450 487524
rect 433333 487459 433399 487460
rect 322197 487388 322263 487389
rect 322197 487384 322244 487388
rect 322308 487386 322314 487388
rect 432137 487386 432203 487389
rect 432270 487386 432276 487388
rect 322197 487328 322202 487384
rect 322197 487324 322244 487328
rect 322308 487326 322354 487386
rect 432137 487384 432276 487386
rect 432137 487328 432142 487384
rect 432198 487328 432276 487384
rect 432137 487326 432276 487328
rect 322308 487324 322314 487326
rect 322197 487323 322263 487324
rect 432137 487323 432203 487326
rect 432270 487324 432276 487326
rect 432340 487324 432346 487388
rect 434713 487386 434779 487389
rect 434846 487386 434852 487388
rect 434713 487384 434852 487386
rect 434713 487328 434718 487384
rect 434774 487328 434852 487384
rect 434713 487326 434852 487328
rect 434713 487323 434779 487326
rect 434846 487324 434852 487326
rect 434916 487324 434922 487388
rect 115606 487188 115612 487252
rect 115676 487250 115682 487252
rect 115841 487250 115907 487253
rect 115676 487248 115907 487250
rect 115676 487192 115846 487248
rect 115902 487192 115907 487248
rect 115676 487190 115907 487192
rect 115676 487188 115682 487190
rect 115841 487187 115907 487190
rect 120574 487188 120580 487252
rect 120644 487250 120650 487252
rect 121361 487250 121427 487253
rect 120644 487248 121427 487250
rect 120644 487192 121366 487248
rect 121422 487192 121427 487248
rect 120644 487190 121427 487192
rect 120644 487188 120650 487190
rect 121361 487187 121427 487190
rect 125542 487188 125548 487252
rect 125612 487250 125618 487252
rect 126881 487250 126947 487253
rect 125612 487248 126947 487250
rect 125612 487192 126886 487248
rect 126942 487192 126947 487248
rect 125612 487190 126947 487192
rect 125612 487188 125618 487190
rect 126881 487187 126947 487190
rect 130510 487188 130516 487252
rect 130580 487250 130586 487252
rect 131021 487250 131087 487253
rect 130580 487248 131087 487250
rect 130580 487192 131026 487248
rect 131082 487192 131087 487248
rect 130580 487190 131087 487192
rect 130580 487188 130586 487190
rect 131021 487187 131087 487190
rect 135478 487188 135484 487252
rect 135548 487250 135554 487252
rect 136541 487250 136607 487253
rect 140681 487252 140747 487253
rect 140630 487250 140636 487252
rect 135548 487248 136607 487250
rect 135548 487192 136546 487248
rect 136602 487192 136607 487248
rect 135548 487190 136607 487192
rect 140590 487190 140636 487250
rect 140700 487248 140747 487252
rect 140742 487192 140747 487248
rect 135548 487188 135554 487190
rect 136541 487187 136607 487190
rect 140630 487188 140636 487190
rect 140700 487188 140747 487192
rect 203006 487188 203012 487252
rect 203076 487250 203082 487252
rect 203517 487250 203583 487253
rect 203076 487248 203583 487250
rect 203076 487192 203522 487248
rect 203578 487192 203583 487248
rect 203076 487190 203583 487192
rect 203076 487188 203082 487190
rect 140681 487187 140747 487188
rect 203517 487187 203583 487190
rect 204897 487250 204963 487253
rect 207657 487252 207723 487253
rect 205398 487250 205404 487252
rect 204897 487248 205404 487250
rect 204897 487192 204902 487248
rect 204958 487192 205404 487248
rect 204897 487190 205404 487192
rect 204897 487187 204963 487190
rect 205398 487188 205404 487190
rect 205468 487188 205474 487252
rect 207606 487250 207612 487252
rect 207566 487190 207612 487250
rect 207676 487248 207723 487252
rect 207718 487192 207723 487248
rect 207606 487188 207612 487190
rect 207676 487188 207723 487192
rect 209998 487188 210004 487252
rect 210068 487250 210074 487252
rect 210417 487250 210483 487253
rect 210068 487248 210483 487250
rect 210068 487192 210422 487248
rect 210478 487192 210483 487248
rect 210068 487190 210483 487192
rect 210068 487188 210074 487190
rect 207657 487187 207723 487188
rect 210417 487187 210483 487190
rect 215334 487188 215340 487252
rect 215404 487250 215410 487252
rect 216581 487250 216647 487253
rect 215404 487248 216647 487250
rect 215404 487192 216586 487248
rect 216642 487192 216647 487248
rect 215404 487190 216647 487192
rect 215404 487188 215410 487190
rect 216581 487187 216647 487190
rect 220486 487188 220492 487252
rect 220556 487250 220562 487252
rect 220721 487250 220787 487253
rect 220556 487248 220787 487250
rect 220556 487192 220726 487248
rect 220782 487192 220787 487248
rect 220556 487190 220787 487192
rect 220556 487188 220562 487190
rect 220721 487187 220787 487190
rect 225454 487188 225460 487252
rect 225524 487250 225530 487252
rect 226241 487250 226307 487253
rect 225524 487248 226307 487250
rect 225524 487192 226246 487248
rect 226302 487192 226307 487248
rect 225524 487190 226307 487192
rect 225524 487188 225530 487190
rect 226241 487187 226307 487190
rect 230606 487188 230612 487252
rect 230676 487250 230682 487252
rect 231761 487250 231827 487253
rect 230676 487248 231827 487250
rect 230676 487192 231766 487248
rect 231822 487192 231827 487248
rect 230676 487190 231827 487192
rect 230676 487188 230682 487190
rect 231761 487187 231827 487190
rect 235574 487188 235580 487252
rect 235644 487250 235650 487252
rect 235901 487250 235967 487253
rect 235644 487248 235967 487250
rect 235644 487192 235906 487248
rect 235962 487192 235967 487248
rect 235644 487190 235967 487192
rect 235644 487188 235650 487190
rect 235901 487187 235967 487190
rect 240542 487188 240548 487252
rect 240612 487250 240618 487252
rect 241421 487250 241487 487253
rect 240612 487248 241487 487250
rect 240612 487192 241426 487248
rect 241482 487192 241487 487248
rect 240612 487190 241487 487192
rect 240612 487188 240618 487190
rect 241421 487187 241487 487190
rect 244641 487250 244707 487253
rect 245510 487250 245516 487252
rect 244641 487248 245516 487250
rect 244641 487192 244646 487248
rect 244702 487192 245516 487248
rect 244641 487190 245516 487192
rect 244641 487187 244707 487190
rect 245510 487188 245516 487190
rect 245580 487188 245586 487252
rect 249793 487250 249859 487253
rect 250478 487250 250484 487252
rect 249793 487248 250484 487250
rect 249793 487192 249798 487248
rect 249854 487192 250484 487248
rect 249793 487190 250484 487192
rect 249793 487187 249859 487190
rect 250478 487188 250484 487190
rect 250548 487188 250554 487252
rect 317638 487188 317644 487252
rect 317708 487250 317714 487252
rect 318057 487250 318123 487253
rect 317708 487248 318123 487250
rect 317708 487192 318062 487248
rect 318118 487192 318123 487248
rect 317708 487190 318123 487192
rect 317708 487188 317714 487190
rect 318057 487187 318123 487190
rect 318926 487188 318932 487252
rect 318996 487250 319002 487252
rect 319437 487250 319503 487253
rect 318996 487248 319503 487250
rect 318996 487192 319442 487248
rect 319498 487192 319503 487248
rect 318996 487190 319503 487192
rect 318996 487188 319002 487190
rect 319437 487187 319503 487190
rect 320817 487250 320883 487253
rect 321134 487250 321140 487252
rect 320817 487248 321140 487250
rect 320817 487192 320822 487248
rect 320878 487192 321140 487248
rect 320817 487190 321140 487192
rect 320817 487187 320883 487190
rect 321134 487188 321140 487190
rect 321204 487188 321210 487252
rect 324313 487250 324379 487253
rect 325182 487250 325188 487252
rect 324313 487248 325188 487250
rect 324313 487192 324318 487248
rect 324374 487192 325188 487248
rect 324313 487190 325188 487192
rect 324313 487187 324379 487190
rect 325182 487188 325188 487190
rect 325252 487188 325258 487252
rect 329833 487250 329899 487253
rect 330518 487250 330524 487252
rect 329833 487248 330524 487250
rect 329833 487192 329838 487248
rect 329894 487192 330524 487248
rect 329833 487190 330524 487192
rect 329833 487187 329899 487190
rect 330518 487188 330524 487190
rect 330588 487188 330594 487252
rect 335353 487250 335419 487253
rect 335486 487250 335492 487252
rect 335353 487248 335492 487250
rect 335353 487192 335358 487248
rect 335414 487192 335492 487248
rect 335353 487190 335492 487192
rect 335353 487187 335419 487190
rect 335486 487188 335492 487190
rect 335556 487188 335562 487252
rect 339493 487250 339559 487253
rect 340454 487250 340460 487252
rect 339493 487248 340460 487250
rect 339493 487192 339498 487248
rect 339554 487192 340460 487248
rect 339493 487190 340460 487192
rect 339493 487187 339559 487190
rect 340454 487188 340460 487190
rect 340524 487188 340530 487252
rect 345013 487250 345079 487253
rect 345606 487250 345612 487252
rect 345013 487248 345612 487250
rect 345013 487192 345018 487248
rect 345074 487192 345612 487248
rect 345013 487190 345612 487192
rect 345013 487187 345079 487190
rect 345606 487188 345612 487190
rect 345676 487188 345682 487252
rect 349153 487250 349219 487253
rect 350390 487250 350396 487252
rect 349153 487248 350396 487250
rect 349153 487192 349158 487248
rect 349214 487192 350396 487248
rect 349153 487190 350396 487192
rect 349153 487187 349219 487190
rect 350390 487188 350396 487190
rect 350460 487188 350466 487252
rect 354673 487250 354739 487253
rect 355542 487250 355548 487252
rect 354673 487248 355548 487250
rect 354673 487192 354678 487248
rect 354734 487192 355548 487248
rect 354673 487190 355548 487192
rect 354673 487187 354739 487190
rect 355542 487188 355548 487190
rect 355612 487188 355618 487252
rect 360193 487250 360259 487253
rect 360510 487250 360516 487252
rect 360193 487248 360516 487250
rect 360193 487192 360198 487248
rect 360254 487192 360516 487248
rect 360193 487190 360516 487192
rect 360193 487187 360259 487190
rect 360510 487188 360516 487190
rect 360580 487188 360586 487252
rect 434713 487250 434779 487253
rect 435214 487250 435220 487252
rect 434713 487248 435220 487250
rect 434713 487192 434718 487248
rect 434774 487192 435220 487248
rect 434713 487190 435220 487192
rect 434713 487187 434779 487190
rect 435214 487188 435220 487190
rect 435284 487188 435290 487252
rect 440233 487250 440299 487253
rect 440366 487250 440372 487252
rect 440233 487248 440372 487250
rect 440233 487192 440238 487248
rect 440294 487192 440372 487248
rect 440233 487190 440372 487192
rect 440233 487187 440299 487190
rect 440366 487188 440372 487190
rect 440436 487188 440442 487252
rect 444373 487250 444439 487253
rect 445518 487250 445524 487252
rect 444373 487248 445524 487250
rect 444373 487192 444378 487248
rect 444434 487192 445524 487248
rect 444373 487190 445524 487192
rect 444373 487187 444439 487190
rect 445518 487188 445524 487190
rect 445588 487188 445594 487252
rect 449893 487250 449959 487253
rect 455413 487252 455479 487253
rect 450486 487250 450492 487252
rect 449893 487248 450492 487250
rect 449893 487192 449898 487248
rect 449954 487192 450492 487248
rect 449893 487190 450492 487192
rect 449893 487187 449959 487190
rect 450486 487188 450492 487190
rect 450556 487188 450562 487252
rect 455413 487250 455460 487252
rect 455368 487248 455460 487250
rect 455368 487192 455418 487248
rect 455368 487190 455460 487192
rect 455413 487188 455460 487190
rect 455524 487188 455530 487252
rect 459553 487250 459619 487253
rect 460422 487250 460428 487252
rect 459553 487248 460428 487250
rect 459553 487192 459558 487248
rect 459614 487192 460428 487248
rect 459553 487190 460428 487192
rect 455413 487187 455479 487188
rect 459553 487187 459619 487190
rect 460422 487188 460428 487190
rect 460492 487188 460498 487252
rect 470593 487250 470659 487253
rect 470726 487250 470732 487252
rect 470593 487248 470732 487250
rect 470593 487192 470598 487248
rect 470654 487192 470732 487248
rect 470593 487190 470732 487192
rect 470593 487187 470659 487190
rect 470726 487188 470732 487190
rect 470796 487188 470802 487252
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2865 462634 2931 462637
rect -960 462632 2931 462634
rect -960 462576 2870 462632
rect 2926 462576 2931 462632
rect -960 462574 2931 462576
rect -960 462484 480 462574
rect 2865 462571 2931 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 232037 454338 232103 454341
rect 382222 454338 382228 454340
rect 232037 454336 382228 454338
rect 232037 454280 232042 454336
rect 232098 454280 382228 454336
rect 232037 454278 382228 454280
rect 232037 454275 232103 454278
rect 382222 454276 382228 454278
rect 382292 454276 382298 454340
rect 232129 454202 232195 454205
rect 382406 454202 382412 454204
rect 232129 454200 382412 454202
rect 232129 454144 232134 454200
rect 232190 454144 382412 454200
rect 232129 454142 382412 454144
rect 232129 454139 232195 454142
rect 382406 454140 382412 454142
rect 382476 454140 382482 454204
rect 225689 454066 225755 454069
rect 383929 454066 383995 454069
rect 225689 454064 383995 454066
rect 225689 454008 225694 454064
rect 225750 454008 383934 454064
rect 383990 454008 383995 454064
rect 225689 454006 383995 454008
rect 225689 454003 225755 454006
rect 383929 454003 383995 454006
rect 297633 452434 297699 452437
rect 297633 452432 300196 452434
rect 297633 452376 297638 452432
rect 297694 452376 300196 452432
rect 297633 452374 300196 452376
rect 297633 452371 297699 452374
rect 384021 452298 384087 452301
rect 383886 452296 384087 452298
rect 383886 452240 384026 452296
rect 384082 452240 384087 452296
rect 383886 452238 384087 452240
rect 383886 451724 383946 452238
rect 384021 452235 384087 452238
rect 234061 449850 234127 449853
rect 297909 449850 297975 449853
rect 234061 449848 297975 449850
rect 234061 449792 234066 449848
rect 234122 449792 297914 449848
rect 297970 449792 297975 449848
rect 234061 449790 297975 449792
rect 234061 449787 234127 449790
rect 297909 449787 297975 449790
rect 255405 449714 255471 449717
rect 256417 449714 256483 449717
rect 292021 449714 292087 449717
rect 255405 449712 292087 449714
rect -960 449578 480 449668
rect 255405 449656 255410 449712
rect 255466 449656 256422 449712
rect 256478 449656 292026 449712
rect 292082 449656 292087 449712
rect 255405 449654 292087 449656
rect 255405 449651 255471 449654
rect 256417 449651 256483 449654
rect 292021 449651 292087 449654
rect 3233 449578 3299 449581
rect -960 449576 3299 449578
rect -960 449520 3238 449576
rect 3294 449520 3299 449576
rect -960 449518 3299 449520
rect -960 449428 480 449518
rect 3233 449515 3299 449518
rect 231669 448762 231735 448765
rect 293166 448762 293172 448764
rect 231669 448760 293172 448762
rect 231669 448704 231674 448760
rect 231730 448704 293172 448760
rect 231669 448702 293172 448704
rect 231669 448699 231735 448702
rect 293166 448700 293172 448702
rect 293236 448700 293242 448764
rect 224401 448626 224467 448629
rect 299381 448626 299447 448629
rect 224401 448624 299447 448626
rect 224401 448568 224406 448624
rect 224462 448568 299386 448624
rect 299442 448568 299447 448624
rect 224401 448566 299447 448568
rect 224401 448563 224467 448566
rect 299381 448563 299447 448566
rect 298001 448354 298067 448357
rect 298001 448352 300196 448354
rect 298001 448296 298006 448352
rect 298062 448296 300196 448352
rect 298001 448294 300196 448296
rect 298001 448291 298067 448294
rect 384021 448218 384087 448221
rect 383886 448216 384087 448218
rect 383886 448160 384026 448216
rect 384082 448160 384087 448216
rect 383886 448158 384087 448160
rect 383886 447644 383946 448158
rect 384021 448155 384087 448158
rect 211153 447266 211219 447269
rect 295977 447266 296043 447269
rect 211153 447264 296043 447266
rect 211153 447208 211158 447264
rect 211214 447208 295982 447264
rect 296038 447208 296043 447264
rect 211153 447206 296043 447208
rect 211153 447203 211219 447206
rect 295977 447203 296043 447206
rect 3366 446660 3372 446724
rect 3436 446722 3442 446724
rect 229737 446722 229803 446725
rect 3436 446720 229803 446722
rect 3436 446664 229742 446720
rect 229798 446664 229803 446720
rect 3436 446662 229803 446664
rect 3436 446660 3442 446662
rect 229737 446659 229803 446662
rect 223297 446586 223363 446589
rect 258574 446586 258580 446588
rect 223297 446584 258580 446586
rect 223297 446528 223302 446584
rect 223358 446528 258580 446584
rect 223297 446526 258580 446528
rect 223297 446523 223363 446526
rect 258574 446524 258580 446526
rect 258644 446524 258650 446588
rect 3509 446450 3575 446453
rect 229185 446450 229251 446453
rect 3509 446448 229251 446450
rect 3509 446392 3514 446448
rect 3570 446392 229190 446448
rect 229246 446392 229251 446448
rect 3509 446390 229251 446392
rect 3509 446387 3575 446390
rect 229185 446387 229251 446390
rect 255497 446450 255563 446453
rect 282126 446450 282132 446452
rect 255497 446448 282132 446450
rect 255497 446392 255502 446448
rect 255558 446392 282132 446448
rect 255497 446390 282132 446392
rect 255497 446387 255563 446390
rect 282126 446388 282132 446390
rect 282196 446388 282202 446452
rect 210417 446314 210483 446317
rect 298829 446314 298895 446317
rect 210417 446312 298895 446314
rect 210417 446256 210422 446312
rect 210478 446256 298834 446312
rect 298890 446256 298895 446312
rect 210417 446254 298895 446256
rect 210417 446251 210483 446254
rect 298829 446251 298895 446254
rect 209129 446178 209195 446181
rect 298502 446178 298508 446180
rect 209129 446176 298508 446178
rect 209129 446120 209134 446176
rect 209190 446120 298508 446176
rect 209129 446118 298508 446120
rect 209129 446115 209195 446118
rect 298502 446116 298508 446118
rect 298572 446116 298578 446180
rect 79317 446042 79383 446045
rect 229369 446042 229435 446045
rect 79317 446040 229435 446042
rect 79317 445984 79322 446040
rect 79378 445984 229374 446040
rect 229430 445984 229435 446040
rect 79317 445982 229435 445984
rect 79317 445979 79383 445982
rect 229369 445979 229435 445982
rect 226241 445906 226307 445909
rect 264094 445906 264100 445908
rect 226241 445904 264100 445906
rect 226241 445848 226246 445904
rect 226302 445848 264100 445904
rect 226241 445846 264100 445848
rect 226241 445843 226307 445846
rect 264094 445844 264100 445846
rect 264164 445844 264170 445908
rect 256785 445770 256851 445773
rect 262622 445770 262628 445772
rect 256785 445768 262628 445770
rect 256785 445712 256790 445768
rect 256846 445712 262628 445768
rect 256785 445710 262628 445712
rect 256785 445707 256851 445710
rect 262622 445708 262628 445710
rect 262692 445708 262698 445772
rect 210049 444954 210115 444957
rect 273897 444954 273963 444957
rect 210049 444952 273963 444954
rect 210049 444896 210054 444952
rect 210110 444896 273902 444952
rect 273958 444896 273963 444952
rect 210049 444894 273963 444896
rect 210049 444891 210115 444894
rect 273897 444891 273963 444894
rect 209681 444818 209747 444821
rect 262438 444818 262444 444820
rect 209681 444816 262444 444818
rect 209681 444760 209686 444816
rect 209742 444760 262444 444816
rect 209681 444758 262444 444760
rect 209681 444755 209747 444758
rect 262438 444756 262444 444758
rect 262508 444756 262514 444820
rect 210233 444682 210299 444685
rect 265617 444682 265683 444685
rect 210233 444680 265683 444682
rect 210233 444624 210238 444680
rect 210294 444624 265622 444680
rect 265678 444624 265683 444680
rect 583520 444668 584960 444908
rect 210233 444622 265683 444624
rect 210233 444619 210299 444622
rect 265617 444619 265683 444622
rect 210785 444546 210851 444549
rect 268377 444546 268443 444549
rect 210785 444544 268443 444546
rect 210785 444488 210790 444544
rect 210846 444488 268382 444544
rect 268438 444488 268443 444544
rect 210785 444486 268443 444488
rect 210785 444483 210851 444486
rect 268377 444483 268443 444486
rect 254393 444410 254459 444413
rect 261518 444410 261524 444412
rect 254393 444408 261524 444410
rect 254393 444352 254398 444408
rect 254454 444352 261524 444408
rect 254393 444350 261524 444352
rect 254393 444347 254459 444350
rect 261518 444348 261524 444350
rect 261588 444348 261594 444412
rect 253473 444274 253539 444277
rect 260046 444274 260052 444276
rect 253473 444272 260052 444274
rect 253473 444216 253478 444272
rect 253534 444216 260052 444272
rect 253473 444214 260052 444216
rect 253473 444211 253539 444214
rect 260046 444212 260052 444214
rect 260116 444212 260122 444276
rect 209497 444138 209563 444141
rect 209630 444138 209636 444140
rect 209497 444136 209636 444138
rect 209497 444080 209502 444136
rect 209558 444080 209636 444136
rect 209497 444078 209636 444080
rect 209497 444075 209563 444078
rect 209630 444076 209636 444078
rect 209700 444076 209706 444140
rect 210601 444138 210667 444141
rect 210734 444138 210740 444140
rect 210601 444136 210740 444138
rect 210601 444080 210606 444136
rect 210662 444080 210740 444136
rect 210601 444078 210740 444080
rect 210601 444075 210667 444078
rect 210734 444076 210740 444078
rect 210804 444076 210810 444140
rect 225505 444138 225571 444141
rect 226701 444138 226767 444141
rect 225505 444136 226767 444138
rect 225505 444080 225510 444136
rect 225566 444080 226706 444136
rect 226762 444080 226767 444136
rect 225505 444078 226767 444080
rect 225505 444075 225571 444078
rect 226701 444075 226767 444078
rect 238017 444138 238083 444141
rect 256417 444140 256483 444141
rect 238150 444138 238156 444140
rect 238017 444136 238156 444138
rect 238017 444080 238022 444136
rect 238078 444080 238156 444136
rect 238017 444078 238156 444080
rect 238017 444075 238083 444078
rect 238150 444076 238156 444078
rect 238220 444076 238226 444140
rect 256366 444138 256372 444140
rect 256326 444078 256372 444138
rect 256436 444136 256483 444140
rect 256478 444080 256483 444136
rect 256366 444076 256372 444078
rect 256436 444076 256483 444080
rect 256417 444075 256483 444076
rect 245469 444004 245535 444005
rect 250989 444004 251055 444005
rect 245469 444000 245516 444004
rect 245580 444002 245586 444004
rect 245469 443944 245474 444000
rect 245469 443940 245516 443944
rect 245580 443942 245626 444002
rect 250989 444000 251036 444004
rect 251100 444002 251106 444004
rect 250989 443944 250994 444000
rect 245580 443940 245586 443942
rect 250989 443940 251036 443944
rect 251100 443942 251146 444002
rect 251100 443940 251106 443942
rect 245469 443939 245535 443940
rect 250989 443939 251055 443940
rect 209405 443866 209471 443869
rect 298737 443866 298803 443869
rect 209405 443864 298803 443866
rect 209405 443808 209410 443864
rect 209466 443808 298742 443864
rect 298798 443808 298803 443864
rect 209405 443806 298803 443808
rect 209405 443803 209471 443806
rect 298737 443803 298803 443806
rect 220118 443668 220124 443732
rect 220188 443730 220194 443732
rect 226333 443730 226399 443733
rect 220188 443728 226399 443730
rect 220188 443672 226338 443728
rect 226394 443672 226399 443728
rect 220188 443670 226399 443672
rect 220188 443668 220194 443670
rect 226333 443667 226399 443670
rect 226701 443730 226767 443733
rect 265801 443730 265867 443733
rect 226701 443728 265867 443730
rect 226701 443672 226706 443728
rect 226762 443672 265806 443728
rect 265862 443672 265867 443728
rect 226701 443670 265867 443672
rect 226701 443667 226767 443670
rect 265801 443667 265867 443670
rect 209957 443594 210023 443597
rect 261334 443594 261340 443596
rect 209957 443592 261340 443594
rect 209957 443536 209962 443592
rect 210018 443536 261340 443592
rect 209957 443534 261340 443536
rect 209957 443531 210023 443534
rect 261334 443532 261340 443534
rect 261404 443532 261410 443596
rect 298001 443594 298067 443597
rect 298001 443592 300196 443594
rect 298001 443536 298006 443592
rect 298062 443536 300196 443592
rect 298001 443534 300196 443536
rect 298001 443531 298067 443534
rect 211061 443458 211127 443461
rect 212349 443458 212415 443461
rect 213637 443458 213703 443461
rect 299289 443458 299355 443461
rect 211061 443456 212274 443458
rect 211061 443400 211066 443456
rect 211122 443400 212274 443456
rect 211061 443398 212274 443400
rect 211061 443395 211127 443398
rect 212214 443186 212274 443398
rect 212349 443456 213562 443458
rect 212349 443400 212354 443456
rect 212410 443400 213562 443456
rect 212349 443398 213562 443400
rect 212349 443395 212415 443398
rect 213502 443322 213562 443398
rect 213637 443456 299355 443458
rect 213637 443400 213642 443456
rect 213698 443400 299294 443456
rect 299350 443400 299355 443456
rect 213637 443398 299355 443400
rect 213637 443395 213703 443398
rect 299289 443395 299355 443398
rect 299105 443322 299171 443325
rect 213502 443320 299171 443322
rect 213502 443264 299110 443320
rect 299166 443264 299171 443320
rect 213502 443262 299171 443264
rect 299105 443259 299171 443262
rect 298921 443186 298987 443189
rect 212214 443184 298987 443186
rect 212214 443128 298926 443184
rect 298982 443128 298987 443184
rect 212214 443126 298987 443128
rect 298921 443123 298987 443126
rect 203374 442988 203380 443052
rect 203444 443050 203450 443052
rect 220118 443050 220124 443052
rect 203444 442990 220124 443050
rect 203444 442988 203450 442990
rect 220118 442988 220124 442990
rect 220188 442988 220194 443052
rect 385309 442914 385375 442917
rect 383916 442912 385375 442914
rect 383916 442856 385314 442912
rect 385370 442856 385375 442912
rect 383916 442854 385375 442856
rect 385309 442851 385375 442854
rect 251030 442716 251036 442780
rect 251100 442778 251106 442780
rect 293125 442778 293191 442781
rect 251100 442776 293191 442778
rect 251100 442720 293130 442776
rect 293186 442720 293191 442776
rect 251100 442718 293191 442720
rect 251100 442716 251106 442718
rect 293125 442715 293191 442718
rect 245510 442580 245516 442644
rect 245580 442642 245586 442644
rect 293769 442642 293835 442645
rect 245580 442640 293835 442642
rect 245580 442584 293774 442640
rect 293830 442584 293835 442640
rect 245580 442582 293835 442584
rect 245580 442580 245586 442582
rect 293769 442579 293835 442582
rect 238150 442444 238156 442508
rect 238220 442506 238226 442508
rect 292941 442506 293007 442509
rect 238220 442504 293007 442506
rect 238220 442448 292946 442504
rect 293002 442448 293007 442504
rect 238220 442446 293007 442448
rect 238220 442444 238226 442446
rect 292941 442443 293007 442446
rect 210734 442308 210740 442372
rect 210804 442370 210810 442372
rect 296069 442370 296135 442373
rect 210804 442368 296135 442370
rect 210804 442312 296074 442368
rect 296130 442312 296135 442368
rect 210804 442310 296135 442312
rect 210804 442308 210810 442310
rect 296069 442307 296135 442310
rect 209630 442172 209636 442236
rect 209700 442234 209706 442236
rect 295926 442234 295932 442236
rect 209700 442174 295932 442234
rect 209700 442172 209706 442174
rect 295926 442172 295932 442174
rect 295996 442172 296002 442236
rect 256366 441628 256372 441692
rect 256436 441690 256442 441692
rect 260230 441690 260236 441692
rect 256436 441630 260236 441690
rect 256436 441628 256442 441630
rect 260230 441628 260236 441630
rect 260300 441628 260306 441692
rect 296805 439514 296871 439517
rect 296805 439512 300196 439514
rect 296805 439456 296810 439512
rect 296866 439456 300196 439512
rect 296805 439454 300196 439456
rect 296805 439451 296871 439454
rect 383886 438701 383946 438804
rect 383886 438696 383995 438701
rect 383886 438640 383934 438696
rect 383990 438640 383995 438696
rect 383886 438638 383995 438640
rect 383929 438635 383995 438638
rect -960 436508 480 436748
rect 296897 434754 296963 434757
rect 296897 434752 300196 434754
rect 296897 434696 296902 434752
rect 296958 434696 300196 434752
rect 296897 434694 300196 434696
rect 296897 434691 296963 434694
rect 385217 434074 385283 434077
rect 383916 434072 385283 434074
rect 383916 434016 385222 434072
rect 385278 434016 385283 434072
rect 383916 434014 385283 434016
rect 385217 434011 385283 434014
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 298001 430674 298067 430677
rect 298001 430672 300196 430674
rect 298001 430616 298006 430672
rect 298062 430616 300196 430672
rect 298001 430614 300196 430616
rect 298001 430611 298067 430614
rect 385125 429994 385191 429997
rect 383916 429992 385191 429994
rect 383916 429936 385130 429992
rect 385186 429936 385191 429992
rect 383916 429934 385191 429936
rect 385125 429931 385191 429934
rect 298001 425914 298067 425917
rect 298001 425912 300196 425914
rect 298001 425856 298006 425912
rect 298062 425856 300196 425912
rect 298001 425854 300196 425856
rect 298001 425851 298067 425854
rect 383326 425716 383332 425780
rect 383396 425716 383402 425780
rect 383334 425204 383394 425716
rect -960 423602 480 423692
rect 3233 423602 3299 423605
rect -960 423600 3299 423602
rect -960 423544 3238 423600
rect 3294 423544 3299 423600
rect -960 423542 3299 423544
rect -960 423452 480 423542
rect 3233 423539 3299 423542
rect 297633 421834 297699 421837
rect 297633 421832 300196 421834
rect 297633 421776 297638 421832
rect 297694 421776 300196 421832
rect 297633 421774 300196 421776
rect 297633 421771 297699 421774
rect 383929 421698 383995 421701
rect 383886 421696 383995 421698
rect 383886 421640 383934 421696
rect 383990 421640 383995 421696
rect 383886 421635 383995 421640
rect 383886 421124 383946 421635
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 297541 417074 297607 417077
rect 297541 417072 300196 417074
rect 297541 417016 297546 417072
rect 297602 417016 300196 417072
rect 297541 417014 300196 417016
rect 297541 417011 297607 417014
rect 385033 416394 385099 416397
rect 383916 416392 385099 416394
rect 383916 416336 385038 416392
rect 385094 416336 385099 416392
rect 383916 416334 385099 416336
rect 385033 416331 385099 416334
rect 297449 412994 297515 412997
rect 297449 412992 300196 412994
rect 297449 412936 297454 412992
rect 297510 412936 300196 412992
rect 297449 412934 300196 412936
rect 297449 412931 297515 412934
rect 383326 412524 383332 412588
rect 383396 412524 383402 412588
rect 383334 412284 383394 412524
rect -960 410546 480 410636
rect 2773 410546 2839 410549
rect -960 410544 2839 410546
rect -960 410488 2778 410544
rect 2834 410488 2839 410544
rect -960 410486 2839 410488
rect -960 410396 480 410486
rect 2773 410483 2839 410486
rect 297357 408234 297423 408237
rect 297357 408232 300196 408234
rect 297357 408176 297362 408232
rect 297418 408176 300196 408232
rect 297357 408174 300196 408176
rect 297357 408171 297423 408174
rect 385033 407554 385099 407557
rect 383916 407552 385099 407554
rect 383916 407496 385038 407552
rect 385094 407496 385099 407552
rect 383916 407494 385099 407496
rect 385033 407491 385099 407494
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect 298001 404154 298067 404157
rect 298001 404152 300196 404154
rect 298001 404096 298006 404152
rect 298062 404096 300196 404152
rect 298001 404094 300196 404096
rect 298001 404091 298067 404094
rect 383334 402932 383394 403444
rect 383326 402868 383332 402932
rect 383396 402868 383402 402932
rect 260046 401508 260052 401572
rect 260116 401570 260122 401572
rect 383326 401570 383332 401572
rect 260116 401510 383332 401570
rect 260116 401508 260122 401510
rect 383326 401508 383332 401510
rect 383396 401508 383402 401572
rect 293125 400890 293191 400893
rect 293125 400888 374010 400890
rect 293125 400832 293130 400888
rect 293186 400832 374010 400888
rect 293125 400830 374010 400832
rect 293125 400827 293191 400830
rect 373950 400754 374010 400830
rect 382733 400754 382799 400757
rect 373950 400752 382799 400754
rect 373950 400696 382738 400752
rect 382794 400696 382799 400752
rect 373950 400694 382799 400696
rect 382733 400691 382799 400694
rect 390553 400346 390619 400349
rect 240918 400344 390619 400346
rect 240918 400288 390558 400344
rect 390614 400288 390619 400344
rect 240918 400286 390619 400288
rect 240777 399938 240843 399941
rect 240918 399938 240978 400286
rect 390553 400283 390619 400286
rect 240777 399936 240978 399938
rect 240777 399880 240782 399936
rect 240838 399880 240978 399936
rect 240777 399878 240978 399880
rect 240777 399875 240843 399878
rect 252870 399876 252876 399940
rect 252940 399938 252946 399940
rect 253473 399938 253539 399941
rect 252940 399936 253539 399938
rect 252940 399880 253478 399936
rect 253534 399880 253539 399936
rect 252940 399878 253539 399880
rect 252940 399876 252946 399878
rect 253473 399875 253539 399878
rect 216949 399258 217015 399261
rect 216814 399256 217015 399258
rect 216814 399200 216954 399256
rect 217010 399200 217015 399256
rect 216814 399198 217015 399200
rect 213913 399122 213979 399125
rect 213913 399120 214114 399122
rect 213913 399064 213918 399120
rect 213974 399064 214114 399120
rect 213913 399062 214114 399064
rect 213913 399059 213979 399062
rect 203425 398850 203491 398853
rect 203425 398848 206018 398850
rect 203425 398792 203430 398848
rect 203486 398792 206018 398848
rect 203425 398790 206018 398792
rect 203425 398787 203491 398790
rect 203701 398714 203767 398717
rect 205817 398714 205883 398717
rect 203701 398712 205883 398714
rect 203701 398656 203706 398712
rect 203762 398656 205822 398712
rect 205878 398656 205883 398712
rect 203701 398654 205883 398656
rect 205958 398714 206018 398790
rect 211889 398714 211955 398717
rect 205958 398712 211955 398714
rect 205958 398656 211894 398712
rect 211950 398656 211955 398712
rect 205958 398654 211955 398656
rect 214054 398714 214114 399062
rect 214465 398986 214531 398989
rect 214465 398984 214850 398986
rect 214465 398928 214470 398984
rect 214526 398928 214850 398984
rect 214465 398926 214850 398928
rect 214465 398923 214531 398926
rect 214465 398850 214531 398853
rect 214790 398850 214850 398926
rect 214465 398848 214850 398850
rect 214465 398792 214470 398848
rect 214526 398792 214850 398848
rect 214465 398790 214850 398792
rect 214465 398787 214531 398790
rect 214598 398714 214604 398716
rect 214054 398654 214604 398714
rect 203701 398651 203767 398654
rect 205817 398651 205883 398654
rect 211889 398651 211955 398654
rect 214598 398652 214604 398654
rect 214668 398652 214674 398716
rect 203517 398578 203583 398581
rect 211797 398578 211863 398581
rect 203517 398576 211863 398578
rect 203517 398520 203522 398576
rect 203578 398520 211802 398576
rect 211858 398520 211863 398576
rect 203517 398518 211863 398520
rect 203517 398515 203583 398518
rect 211797 398515 211863 398518
rect 202137 398442 202203 398445
rect 205582 398442 205588 398444
rect 202137 398440 205588 398442
rect 202137 398384 202142 398440
rect 202198 398384 205588 398440
rect 202137 398382 205588 398384
rect 202137 398379 202203 398382
rect 205582 398380 205588 398382
rect 205652 398380 205658 398444
rect 205817 398442 205883 398445
rect 212809 398442 212875 398445
rect 205817 398440 212875 398442
rect 205817 398384 205822 398440
rect 205878 398384 212814 398440
rect 212870 398384 212875 398440
rect 205817 398382 212875 398384
rect 205817 398379 205883 398382
rect 212809 398379 212875 398382
rect 188337 398306 188403 398309
rect 211153 398306 211219 398309
rect 188337 398304 211219 398306
rect 188337 398248 188342 398304
rect 188398 398248 211158 398304
rect 211214 398248 211219 398304
rect 188337 398246 211219 398248
rect 188337 398243 188403 398246
rect 211153 398243 211219 398246
rect 211286 398244 211292 398308
rect 211356 398306 211362 398308
rect 211429 398306 211495 398309
rect 211356 398304 211495 398306
rect 211356 398248 211434 398304
rect 211490 398248 211495 398304
rect 211356 398246 211495 398248
rect 211356 398244 211362 398246
rect 211429 398243 211495 398246
rect 178677 398170 178743 398173
rect 178677 398168 200130 398170
rect 178677 398112 178682 398168
rect 178738 398112 200130 398168
rect 178677 398110 200130 398112
rect 178677 398107 178743 398110
rect 200070 398034 200130 398110
rect 205582 398108 205588 398172
rect 205652 398170 205658 398172
rect 213361 398170 213427 398173
rect 215845 398170 215911 398173
rect 205652 398168 213427 398170
rect 205652 398112 213366 398168
rect 213422 398112 213427 398168
rect 205652 398110 213427 398112
rect 205652 398108 205658 398110
rect 213361 398107 213427 398110
rect 213686 398168 215911 398170
rect 213686 398112 215850 398168
rect 215906 398112 215911 398168
rect 213686 398110 215911 398112
rect 211521 398034 211587 398037
rect 200070 398032 211587 398034
rect 200070 397976 211526 398032
rect 211582 397976 211587 398032
rect 200070 397974 211587 397976
rect 211521 397971 211587 397974
rect 212441 398034 212507 398037
rect 213686 398034 213746 398110
rect 215845 398107 215911 398110
rect 212441 398032 213746 398034
rect 212441 397976 212446 398032
rect 212502 397976 213746 398032
rect 212441 397974 213746 397976
rect 214005 398034 214071 398037
rect 216814 398034 216874 399198
rect 216949 399195 217015 399198
rect 252553 399258 252619 399261
rect 252686 399258 252692 399260
rect 252553 399256 252692 399258
rect 252553 399200 252558 399256
rect 252614 399200 252692 399256
rect 252553 399198 252692 399200
rect 252553 399195 252619 399198
rect 252686 399196 252692 399198
rect 252756 399196 252762 399260
rect 248505 399122 248571 399125
rect 329005 399122 329071 399125
rect 248505 399120 253306 399122
rect 248505 399064 248510 399120
rect 248566 399064 253306 399120
rect 248505 399062 253306 399064
rect 248505 399059 248571 399062
rect 243905 398986 243971 398989
rect 243905 398984 244106 398986
rect 243905 398928 243910 398984
rect 243966 398928 244106 398984
rect 243905 398926 244106 398928
rect 243905 398923 243971 398926
rect 244046 398714 244106 398926
rect 250161 398850 250227 398853
rect 252645 398852 252711 398853
rect 250294 398850 250300 398852
rect 250161 398848 250300 398850
rect 250161 398792 250166 398848
rect 250222 398792 250300 398848
rect 250161 398790 250300 398792
rect 250161 398787 250227 398790
rect 250294 398788 250300 398790
rect 250364 398788 250370 398852
rect 252645 398848 252692 398852
rect 252756 398850 252762 398852
rect 252645 398792 252650 398848
rect 252645 398788 252692 398792
rect 252756 398790 252802 398850
rect 252756 398788 252762 398790
rect 252645 398787 252711 398788
rect 244365 398714 244431 398717
rect 244046 398712 244431 398714
rect 244046 398656 244370 398712
rect 244426 398656 244431 398712
rect 244046 398654 244431 398656
rect 244365 398651 244431 398654
rect 252737 398714 252803 398717
rect 252870 398714 252876 398716
rect 252737 398712 252876 398714
rect 252737 398656 252742 398712
rect 252798 398656 252876 398712
rect 252737 398654 252876 398656
rect 252737 398651 252803 398654
rect 252870 398652 252876 398654
rect 252940 398652 252946 398716
rect 253246 398714 253306 399062
rect 311850 399120 329071 399122
rect 311850 399064 329010 399120
rect 329066 399064 329071 399120
rect 311850 399062 329071 399064
rect 258574 398924 258580 398988
rect 258644 398986 258650 398988
rect 311850 398986 311910 399062
rect 329005 399059 329071 399062
rect 258644 398926 311910 398986
rect 312126 398926 321570 398986
rect 258644 398924 258650 398926
rect 264094 398788 264100 398852
rect 264164 398850 264170 398852
rect 312126 398850 312186 398926
rect 264164 398790 312186 398850
rect 321510 398850 321570 398926
rect 321694 398926 331230 398986
rect 321694 398850 321754 398926
rect 321510 398790 321754 398850
rect 331170 398850 331230 398926
rect 337377 398850 337443 398853
rect 331170 398848 337443 398850
rect 331170 398792 337382 398848
rect 337438 398792 337443 398848
rect 331170 398790 337443 398792
rect 264164 398788 264170 398790
rect 337377 398787 337443 398790
rect 253246 398654 258090 398714
rect 228582 398516 228588 398580
rect 228652 398578 228658 398580
rect 233877 398578 233943 398581
rect 228652 398576 233943 398578
rect 228652 398520 233882 398576
rect 233938 398520 233943 398576
rect 228652 398518 233943 398520
rect 228652 398516 228658 398518
rect 233877 398515 233943 398518
rect 248781 398578 248847 398581
rect 248781 398576 256434 398578
rect 248781 398520 248786 398576
rect 248842 398520 256434 398576
rect 248781 398518 256434 398520
rect 248781 398515 248847 398518
rect 253422 398380 253428 398444
rect 253492 398442 253498 398444
rect 253841 398442 253907 398445
rect 253492 398440 253907 398442
rect 253492 398384 253846 398440
rect 253902 398384 253907 398440
rect 253492 398382 253907 398384
rect 253492 398380 253498 398382
rect 253841 398379 253907 398382
rect 246481 398306 246547 398309
rect 246982 398306 246988 398308
rect 246481 398304 246988 398306
rect 246481 398248 246486 398304
rect 246542 398248 246988 398304
rect 246481 398246 246988 398248
rect 246481 398243 246547 398246
rect 246982 398244 246988 398246
rect 247052 398244 247058 398308
rect 251265 398306 251331 398309
rect 256233 398306 256299 398309
rect 251265 398304 256299 398306
rect 251265 398248 251270 398304
rect 251326 398248 256238 398304
rect 256294 398248 256299 398304
rect 251265 398246 256299 398248
rect 251265 398243 251331 398246
rect 256233 398243 256299 398246
rect 236729 398170 236795 398173
rect 214005 398032 216874 398034
rect 214005 397976 214010 398032
rect 214066 397976 216874 398032
rect 214005 397974 216874 397976
rect 229510 398168 236795 398170
rect 229510 398112 236734 398168
rect 236790 398112 236795 398168
rect 229510 398110 236795 398112
rect 212441 397971 212507 397974
rect 214005 397971 214071 397974
rect 211153 397898 211219 397901
rect 213913 397898 213979 397901
rect 211153 397896 213979 397898
rect 211153 397840 211158 397896
rect 211214 397840 213918 397896
rect 213974 397840 213979 397896
rect 211153 397838 213979 397840
rect 211153 397835 211219 397838
rect 213913 397835 213979 397838
rect 216622 397836 216628 397900
rect 216692 397898 216698 397900
rect 217041 397898 217107 397901
rect 216692 397896 217107 397898
rect 216692 397840 217046 397896
rect 217102 397840 217107 397896
rect 216692 397838 217107 397840
rect 216692 397836 216698 397838
rect 217041 397835 217107 397838
rect 223573 397898 223639 397901
rect 223982 397898 223988 397900
rect 223573 397896 223988 397898
rect 223573 397840 223578 397896
rect 223634 397840 223988 397896
rect 223573 397838 223988 397840
rect 223573 397835 223639 397838
rect 223982 397836 223988 397838
rect 224052 397836 224058 397900
rect 224902 397836 224908 397900
rect 224972 397898 224978 397900
rect 225413 397898 225479 397901
rect 224972 397896 225479 397898
rect 224972 397840 225418 397896
rect 225474 397840 225479 397896
rect 224972 397838 225479 397840
rect 224972 397836 224978 397838
rect 225413 397835 225479 397838
rect 228766 397836 228772 397900
rect 228836 397898 228842 397900
rect 229001 397898 229067 397901
rect 228836 397896 229067 397898
rect 228836 397840 229006 397896
rect 229062 397840 229067 397896
rect 228836 397838 229067 397840
rect 228836 397836 228842 397838
rect 229001 397835 229067 397838
rect 211245 397762 211311 397765
rect 211654 397762 211660 397764
rect 211245 397760 211660 397762
rect 211245 397704 211250 397760
rect 211306 397704 211660 397760
rect 211245 397702 211660 397704
rect 211245 397699 211311 397702
rect 211654 397700 211660 397702
rect 211724 397700 211730 397764
rect 212533 397762 212599 397765
rect 212758 397762 212764 397764
rect 212533 397760 212764 397762
rect 212533 397704 212538 397760
rect 212594 397704 212764 397760
rect 212533 397702 212764 397704
rect 212533 397699 212599 397702
rect 212758 397700 212764 397702
rect 212828 397700 212834 397764
rect 214046 397700 214052 397764
rect 214116 397762 214122 397764
rect 214281 397762 214347 397765
rect 214116 397760 214347 397762
rect 214116 397704 214286 397760
rect 214342 397704 214347 397760
rect 214116 397702 214347 397704
rect 214116 397700 214122 397702
rect 214281 397699 214347 397702
rect 215334 397700 215340 397764
rect 215404 397762 215410 397764
rect 215569 397762 215635 397765
rect 215404 397760 215635 397762
rect 215404 397704 215574 397760
rect 215630 397704 215635 397760
rect 215404 397702 215635 397704
rect 215404 397700 215410 397702
rect 215569 397699 215635 397702
rect 216673 397762 216739 397765
rect 216990 397762 216996 397764
rect 216673 397760 216996 397762
rect 216673 397704 216678 397760
rect 216734 397704 216996 397760
rect 216673 397702 216996 397704
rect 216673 397699 216739 397702
rect 216990 397700 216996 397702
rect 217060 397700 217066 397764
rect 222193 397762 222259 397765
rect 223062 397762 223068 397764
rect 222193 397760 223068 397762
rect 222193 397704 222198 397760
rect 222254 397704 223068 397760
rect 222193 397702 223068 397704
rect 222193 397699 222259 397702
rect 223062 397700 223068 397702
rect 223132 397700 223138 397764
rect 223849 397762 223915 397765
rect 224166 397762 224172 397764
rect 223849 397760 224172 397762
rect 223849 397704 223854 397760
rect 223910 397704 224172 397760
rect 223849 397702 224172 397704
rect 223849 397699 223915 397702
rect 224166 397700 224172 397702
rect 224236 397700 224242 397764
rect 224953 397762 225019 397765
rect 225270 397762 225276 397764
rect 224953 397760 225276 397762
rect 224953 397704 224958 397760
rect 225014 397704 225276 397760
rect 224953 397702 225276 397704
rect 224953 397699 225019 397702
rect 225270 397700 225276 397702
rect 225340 397700 225346 397764
rect 228398 397700 228404 397764
rect 228468 397762 228474 397764
rect 229510 397762 229570 398110
rect 236729 398107 236795 398110
rect 249885 398170 249951 398173
rect 256374 398170 256434 398518
rect 258030 398306 258090 398654
rect 260230 398652 260236 398716
rect 260300 398714 260306 398716
rect 374729 398714 374795 398717
rect 260300 398712 374795 398714
rect 260300 398656 374734 398712
rect 374790 398656 374795 398712
rect 260300 398654 374795 398656
rect 260300 398652 260306 398654
rect 374729 398651 374795 398654
rect 261518 398516 261524 398580
rect 261588 398578 261594 398580
rect 316125 398578 316191 398581
rect 261588 398576 316191 398578
rect 261588 398520 316130 398576
rect 316186 398520 316191 398576
rect 261588 398518 316191 398520
rect 261588 398516 261594 398518
rect 316125 398515 316191 398518
rect 489913 398306 489979 398309
rect 258030 398304 489979 398306
rect 258030 398248 489918 398304
rect 489974 398248 489979 398304
rect 258030 398246 489979 398248
rect 489913 398243 489979 398246
rect 494053 398170 494119 398173
rect 249885 398168 256250 398170
rect 249885 398112 249890 398168
rect 249946 398112 256250 398168
rect 249885 398110 256250 398112
rect 256374 398168 494119 398170
rect 256374 398112 494058 398168
rect 494114 398112 494119 398168
rect 256374 398110 494119 398112
rect 249885 398107 249951 398110
rect 230197 398034 230263 398037
rect 230422 398034 230428 398036
rect 230197 398032 230428 398034
rect 230197 397976 230202 398032
rect 230258 397976 230428 398032
rect 230197 397974 230428 397976
rect 230197 397971 230263 397974
rect 230422 397972 230428 397974
rect 230492 397972 230498 398036
rect 232957 398034 233023 398037
rect 233182 398034 233188 398036
rect 232957 398032 233188 398034
rect 232957 397976 232962 398032
rect 233018 397976 233188 398032
rect 232957 397974 233188 397976
rect 232957 397971 233023 397974
rect 233182 397972 233188 397974
rect 233252 397972 233258 398036
rect 247953 398034 248019 398037
rect 254025 398034 254091 398037
rect 256049 398034 256115 398037
rect 247953 398032 253950 398034
rect 247953 397976 247958 398032
rect 248014 397976 253950 398032
rect 247953 397974 253950 397976
rect 247953 397971 248019 397974
rect 234705 397898 234771 397901
rect 228468 397702 229570 397762
rect 229694 397896 234771 397898
rect 229694 397840 234710 397896
rect 234766 397840 234771 397896
rect 229694 397838 234771 397840
rect 228468 397700 228474 397702
rect -960 397490 480 397580
rect 209814 397564 209820 397628
rect 209884 397626 209890 397628
rect 210325 397626 210391 397629
rect 209884 397624 210391 397626
rect 209884 397568 210330 397624
rect 210386 397568 210391 397624
rect 209884 397566 210391 397568
rect 209884 397564 209890 397566
rect 210325 397563 210391 397566
rect 211286 397564 211292 397628
rect 211356 397626 211362 397628
rect 211613 397626 211679 397629
rect 211356 397624 211679 397626
rect 211356 397568 211618 397624
rect 211674 397568 211679 397624
rect 211356 397566 211679 397568
rect 211356 397564 211362 397566
rect 211613 397563 211679 397566
rect 211797 397626 211863 397629
rect 212993 397626 213059 397629
rect 214005 397626 214071 397629
rect 211797 397624 213059 397626
rect 211797 397568 211802 397624
rect 211858 397568 212998 397624
rect 213054 397568 213059 397624
rect 211797 397566 213059 397568
rect 211797 397563 211863 397566
rect 212993 397563 213059 397566
rect 213134 397624 214071 397626
rect 213134 397568 214010 397624
rect 214066 397568 214071 397624
rect 213134 397566 214071 397568
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 25497 397490 25563 397493
rect 203425 397490 203491 397493
rect 25497 397488 203491 397490
rect 25497 397432 25502 397488
rect 25558 397432 203430 397488
rect 203486 397432 203491 397488
rect 25497 397430 203491 397432
rect 25497 397427 25563 397430
rect 203425 397427 203491 397430
rect 209998 397428 210004 397492
rect 210068 397490 210074 397492
rect 210417 397490 210483 397493
rect 210068 397488 210483 397490
rect 210068 397432 210422 397488
rect 210478 397432 210483 397488
rect 210068 397430 210483 397432
rect 210068 397428 210074 397430
rect 210417 397427 210483 397430
rect 211337 397490 211403 397493
rect 212625 397492 212691 397493
rect 211470 397490 211476 397492
rect 211337 397488 211476 397490
rect 211337 397432 211342 397488
rect 211398 397432 211476 397488
rect 211337 397430 211476 397432
rect 211337 397427 211403 397430
rect 211470 397428 211476 397430
rect 211540 397428 211546 397492
rect 212574 397490 212580 397492
rect 212534 397430 212580 397490
rect 212644 397488 212691 397492
rect 213134 397490 213194 397566
rect 214005 397563 214071 397566
rect 214189 397626 214255 397629
rect 214414 397626 214420 397628
rect 214189 397624 214420 397626
rect 214189 397568 214194 397624
rect 214250 397568 214420 397624
rect 214189 397566 214420 397568
rect 214189 397563 214255 397566
rect 214414 397564 214420 397566
rect 214484 397564 214490 397628
rect 215477 397626 215543 397629
rect 215702 397626 215708 397628
rect 215477 397624 215708 397626
rect 215477 397568 215482 397624
rect 215538 397568 215708 397624
rect 215477 397566 215708 397568
rect 215477 397563 215543 397566
rect 215702 397564 215708 397566
rect 215772 397564 215778 397628
rect 216857 397626 216923 397629
rect 217174 397626 217180 397628
rect 216857 397624 217180 397626
rect 216857 397568 216862 397624
rect 216918 397568 217180 397624
rect 216857 397566 217180 397568
rect 216857 397563 216923 397566
rect 217174 397564 217180 397566
rect 217244 397564 217250 397628
rect 218237 397626 218303 397629
rect 218830 397626 218836 397628
rect 218237 397624 218836 397626
rect 218237 397568 218242 397624
rect 218298 397568 218836 397624
rect 218237 397566 218836 397568
rect 218237 397563 218303 397566
rect 218830 397564 218836 397566
rect 218900 397564 218906 397628
rect 219566 397564 219572 397628
rect 219636 397626 219642 397628
rect 219801 397626 219867 397629
rect 220905 397628 220971 397629
rect 220854 397626 220860 397628
rect 219636 397624 219867 397626
rect 219636 397568 219806 397624
rect 219862 397568 219867 397624
rect 219636 397566 219867 397568
rect 220814 397566 220860 397626
rect 220924 397624 220971 397628
rect 220966 397568 220971 397624
rect 219636 397564 219642 397566
rect 219801 397563 219867 397566
rect 220854 397564 220860 397566
rect 220924 397564 220971 397568
rect 220905 397563 220971 397564
rect 221089 397626 221155 397629
rect 221406 397626 221412 397628
rect 221089 397624 221412 397626
rect 221089 397568 221094 397624
rect 221150 397568 221412 397624
rect 221089 397566 221412 397568
rect 221089 397563 221155 397566
rect 221406 397564 221412 397566
rect 221476 397564 221482 397628
rect 223614 397564 223620 397628
rect 223684 397626 223690 397628
rect 223941 397626 224007 397629
rect 223684 397624 224007 397626
rect 223684 397568 223946 397624
rect 224002 397568 224007 397624
rect 223684 397566 224007 397568
rect 223684 397564 223690 397566
rect 223941 397563 224007 397566
rect 225229 397626 225295 397629
rect 225454 397626 225460 397628
rect 225229 397624 225460 397626
rect 225229 397568 225234 397624
rect 225290 397568 225460 397624
rect 225229 397566 225460 397568
rect 225229 397563 225295 397566
rect 225454 397564 225460 397566
rect 225524 397564 225530 397628
rect 226558 397564 226564 397628
rect 226628 397626 226634 397628
rect 229694 397626 229754 397838
rect 234705 397835 234771 397838
rect 242382 397836 242388 397900
rect 242452 397898 242458 397900
rect 242801 397898 242867 397901
rect 242452 397896 242867 397898
rect 242452 397840 242806 397896
rect 242862 397840 242867 397896
rect 242452 397838 242867 397840
rect 242452 397836 242458 397838
rect 242801 397835 242867 397838
rect 247718 397836 247724 397900
rect 247788 397898 247794 397900
rect 248321 397898 248387 397901
rect 247788 397896 248387 397898
rect 247788 397840 248326 397896
rect 248382 397840 248387 397896
rect 247788 397838 248387 397840
rect 247788 397836 247794 397838
rect 248321 397835 248387 397838
rect 250478 397836 250484 397900
rect 250548 397898 250554 397900
rect 250897 397898 250963 397901
rect 250548 397896 250963 397898
rect 250548 397840 250902 397896
rect 250958 397840 250963 397896
rect 250548 397838 250963 397840
rect 250548 397836 250554 397838
rect 250897 397835 250963 397838
rect 251766 397836 251772 397900
rect 251836 397898 251842 397900
rect 252185 397898 252251 397901
rect 251836 397896 252251 397898
rect 251836 397840 252190 397896
rect 252246 397840 252251 397896
rect 251836 397838 252251 397840
rect 251836 397836 251842 397838
rect 252185 397835 252251 397838
rect 230054 397700 230060 397764
rect 230124 397762 230130 397764
rect 230381 397762 230447 397765
rect 230124 397760 230447 397762
rect 230124 397704 230386 397760
rect 230442 397704 230447 397760
rect 230124 397702 230447 397704
rect 230124 397700 230130 397702
rect 230381 397699 230447 397702
rect 230606 397700 230612 397764
rect 230676 397762 230682 397764
rect 231577 397762 231643 397765
rect 230676 397760 231643 397762
rect 230676 397704 231582 397760
rect 231638 397704 231643 397760
rect 230676 397702 231643 397704
rect 230676 397700 230682 397702
rect 231577 397699 231643 397702
rect 232814 397700 232820 397764
rect 232884 397762 232890 397764
rect 233141 397762 233207 397765
rect 232884 397760 233207 397762
rect 232884 397704 233146 397760
rect 233202 397704 233207 397760
rect 232884 397702 233207 397704
rect 232884 397700 232890 397702
rect 233141 397699 233207 397702
rect 233918 397700 233924 397764
rect 233988 397762 233994 397764
rect 234429 397762 234495 397765
rect 233988 397760 234495 397762
rect 233988 397704 234434 397760
rect 234490 397704 234495 397760
rect 233988 397702 234495 397704
rect 233988 397700 233994 397702
rect 234429 397699 234495 397702
rect 235206 397700 235212 397764
rect 235276 397762 235282 397764
rect 235901 397762 235967 397765
rect 235276 397760 235967 397762
rect 235276 397704 235906 397760
rect 235962 397704 235967 397760
rect 235276 397702 235967 397704
rect 235276 397700 235282 397702
rect 235901 397699 235967 397702
rect 236862 397700 236868 397764
rect 236932 397762 236938 397764
rect 237097 397762 237163 397765
rect 236932 397760 237163 397762
rect 236932 397704 237102 397760
rect 237158 397704 237163 397760
rect 236932 397702 237163 397704
rect 236932 397700 236938 397702
rect 237097 397699 237163 397702
rect 238150 397700 238156 397764
rect 238220 397762 238226 397764
rect 238385 397762 238451 397765
rect 238220 397760 238451 397762
rect 238220 397704 238390 397760
rect 238446 397704 238451 397760
rect 238220 397702 238451 397704
rect 238220 397700 238226 397702
rect 238385 397699 238451 397702
rect 242198 397700 242204 397764
rect 242268 397762 242274 397764
rect 242525 397762 242591 397765
rect 242268 397760 242591 397762
rect 242268 397704 242530 397760
rect 242586 397704 242591 397760
rect 242268 397702 242591 397704
rect 242268 397700 242274 397702
rect 242525 397699 242591 397702
rect 243670 397700 243676 397764
rect 243740 397762 243746 397764
rect 244181 397762 244247 397765
rect 243740 397760 244247 397762
rect 243740 397704 244186 397760
rect 244242 397704 244247 397760
rect 243740 397702 244247 397704
rect 243740 397700 243746 397702
rect 244181 397699 244247 397702
rect 246430 397700 246436 397764
rect 246500 397762 246506 397764
rect 246941 397762 247007 397765
rect 246500 397760 247007 397762
rect 246500 397704 246946 397760
rect 247002 397704 247007 397760
rect 246500 397702 247007 397704
rect 246500 397700 246506 397702
rect 246941 397699 247007 397702
rect 247902 397700 247908 397764
rect 247972 397762 247978 397764
rect 248137 397762 248203 397765
rect 247972 397760 248203 397762
rect 247972 397704 248142 397760
rect 248198 397704 248203 397760
rect 247972 397702 248203 397704
rect 247972 397700 247978 397702
rect 248137 397699 248203 397702
rect 248638 397700 248644 397764
rect 248708 397762 248714 397764
rect 249701 397762 249767 397765
rect 248708 397760 249767 397762
rect 248708 397704 249706 397760
rect 249762 397704 249767 397760
rect 248708 397702 249767 397704
rect 248708 397700 248714 397702
rect 249701 397699 249767 397702
rect 250662 397700 250668 397764
rect 250732 397762 250738 397764
rect 251081 397762 251147 397765
rect 250732 397760 251147 397762
rect 250732 397704 251086 397760
rect 251142 397704 251147 397760
rect 250732 397702 251147 397704
rect 250732 397700 250738 397702
rect 251081 397699 251147 397702
rect 251950 397700 251956 397764
rect 252020 397762 252026 397764
rect 252277 397762 252343 397765
rect 252020 397760 252343 397762
rect 252020 397704 252282 397760
rect 252338 397704 252343 397760
rect 252020 397702 252343 397704
rect 252020 397700 252026 397702
rect 252277 397699 252343 397702
rect 253238 397700 253244 397764
rect 253308 397762 253314 397764
rect 253749 397762 253815 397765
rect 253308 397760 253815 397762
rect 253308 397704 253754 397760
rect 253810 397704 253815 397760
rect 253308 397702 253815 397704
rect 253308 397700 253314 397702
rect 253749 397699 253815 397702
rect 226628 397566 229754 397626
rect 226628 397564 226634 397566
rect 229870 397564 229876 397628
rect 229940 397626 229946 397628
rect 230105 397626 230171 397629
rect 229940 397624 230171 397626
rect 229940 397568 230110 397624
rect 230166 397568 230171 397624
rect 229940 397566 230171 397568
rect 229940 397564 229946 397566
rect 230105 397563 230171 397566
rect 230790 397564 230796 397628
rect 230860 397626 230866 397628
rect 231761 397626 231827 397629
rect 230860 397624 231827 397626
rect 230860 397568 231766 397624
rect 231822 397568 231827 397624
rect 230860 397566 231827 397568
rect 230860 397564 230866 397566
rect 231761 397563 231827 397566
rect 232630 397564 232636 397628
rect 232700 397626 232706 397628
rect 232865 397626 232931 397629
rect 232700 397624 232931 397626
rect 232700 397568 232870 397624
rect 232926 397568 232931 397624
rect 232700 397566 232931 397568
rect 232700 397564 232706 397566
rect 232865 397563 232931 397566
rect 234102 397564 234108 397628
rect 234172 397626 234178 397628
rect 234337 397626 234403 397629
rect 234172 397624 234403 397626
rect 234172 397568 234342 397624
rect 234398 397568 234403 397624
rect 234172 397566 234403 397568
rect 234172 397564 234178 397566
rect 234337 397563 234403 397566
rect 235390 397564 235396 397628
rect 235460 397626 235466 397628
rect 235717 397626 235783 397629
rect 235460 397624 235783 397626
rect 235460 397568 235722 397624
rect 235778 397568 235783 397624
rect 235460 397566 235783 397568
rect 235460 397564 235466 397566
rect 235717 397563 235783 397566
rect 237046 397564 237052 397628
rect 237116 397626 237122 397628
rect 237281 397626 237347 397629
rect 237116 397624 237347 397626
rect 237116 397568 237286 397624
rect 237342 397568 237347 397624
rect 237116 397566 237347 397568
rect 237116 397564 237122 397566
rect 237281 397563 237347 397566
rect 238334 397564 238340 397628
rect 238404 397626 238410 397628
rect 238477 397626 238543 397629
rect 238404 397624 238543 397626
rect 238404 397568 238482 397624
rect 238538 397568 238543 397624
rect 238404 397566 238543 397568
rect 238404 397564 238410 397566
rect 238477 397563 238543 397566
rect 239806 397564 239812 397628
rect 239876 397626 239882 397628
rect 240041 397626 240107 397629
rect 239876 397624 240107 397626
rect 239876 397568 240046 397624
rect 240102 397568 240107 397624
rect 239876 397566 240107 397568
rect 239876 397564 239882 397566
rect 240041 397563 240107 397566
rect 242433 397626 242499 397629
rect 244089 397628 244155 397629
rect 246665 397628 246731 397629
rect 242750 397626 242756 397628
rect 242433 397624 242756 397626
rect 242433 397568 242438 397624
rect 242494 397568 242756 397624
rect 242433 397566 242756 397568
rect 242433 397563 242499 397566
rect 242750 397564 242756 397566
rect 242820 397564 242826 397628
rect 244038 397626 244044 397628
rect 243998 397566 244044 397626
rect 244108 397624 244155 397628
rect 246614 397626 246620 397628
rect 244150 397568 244155 397624
rect 244038 397564 244044 397566
rect 244108 397564 244155 397568
rect 246574 397566 246620 397626
rect 246684 397624 246731 397628
rect 248045 397628 248111 397629
rect 248045 397626 248092 397628
rect 246726 397568 246731 397624
rect 246614 397564 246620 397566
rect 246684 397564 246731 397568
rect 248000 397624 248092 397626
rect 248000 397568 248050 397624
rect 248000 397566 248092 397568
rect 244089 397563 244155 397564
rect 246665 397563 246731 397564
rect 248045 397564 248092 397566
rect 248156 397564 248162 397628
rect 248822 397564 248828 397628
rect 248892 397626 248898 397628
rect 249517 397626 249583 397629
rect 250805 397628 250871 397629
rect 250805 397626 250852 397628
rect 248892 397624 249583 397626
rect 248892 397568 249522 397624
rect 249578 397568 249583 397624
rect 248892 397566 249583 397568
rect 250760 397624 250852 397626
rect 250760 397568 250810 397624
rect 250760 397566 250852 397568
rect 248892 397564 248898 397566
rect 248045 397563 248111 397564
rect 249517 397563 249583 397566
rect 250805 397564 250852 397566
rect 250916 397564 250922 397628
rect 252134 397564 252140 397628
rect 252204 397626 252210 397628
rect 252461 397626 252527 397629
rect 252204 397624 252527 397626
rect 252204 397568 252466 397624
rect 252522 397568 252527 397624
rect 252204 397566 252527 397568
rect 252204 397564 252210 397566
rect 250805 397563 250871 397564
rect 252461 397563 252527 397566
rect 212686 397432 212691 397488
rect 212574 397428 212580 397430
rect 212644 397428 212691 397432
rect 212625 397427 212691 397428
rect 212766 397430 213194 397490
rect 214097 397490 214163 397493
rect 214230 397490 214236 397492
rect 214097 397488 214236 397490
rect 214097 397432 214102 397488
rect 214158 397432 214236 397488
rect 214097 397430 214236 397432
rect 210417 397354 210483 397357
rect 212766 397354 212826 397430
rect 214097 397427 214163 397430
rect 214230 397428 214236 397430
rect 214300 397428 214306 397492
rect 215293 397490 215359 397493
rect 216765 397492 216831 397493
rect 215518 397490 215524 397492
rect 215293 397488 215524 397490
rect 215293 397432 215298 397488
rect 215354 397432 215524 397488
rect 215293 397430 215524 397432
rect 215293 397427 215359 397430
rect 215518 397428 215524 397430
rect 215588 397428 215594 397492
rect 216765 397490 216812 397492
rect 216720 397488 216812 397490
rect 216720 397432 216770 397488
rect 216720 397430 216812 397432
rect 216765 397428 216812 397430
rect 216876 397428 216882 397492
rect 218053 397490 218119 397493
rect 218646 397490 218652 397492
rect 218053 397488 218652 397490
rect 218053 397432 218058 397488
rect 218114 397432 218652 397488
rect 218053 397430 218652 397432
rect 216765 397427 216831 397428
rect 218053 397427 218119 397430
rect 218646 397428 218652 397430
rect 218716 397428 218722 397492
rect 219382 397428 219388 397492
rect 219452 397490 219458 397492
rect 219525 397490 219591 397493
rect 219709 397492 219775 397493
rect 220997 397492 221063 397493
rect 221181 397492 221247 397493
rect 219709 397490 219756 397492
rect 219452 397488 219591 397490
rect 219452 397432 219530 397488
rect 219586 397432 219591 397488
rect 219452 397430 219591 397432
rect 219664 397488 219756 397490
rect 219664 397432 219714 397488
rect 219664 397430 219756 397432
rect 219452 397428 219458 397430
rect 219525 397427 219591 397430
rect 219709 397428 219756 397430
rect 219820 397428 219826 397492
rect 220997 397490 221044 397492
rect 220952 397488 221044 397490
rect 220952 397432 221002 397488
rect 220952 397430 221044 397432
rect 220997 397428 221044 397430
rect 221108 397428 221114 397492
rect 221181 397488 221228 397492
rect 221292 397490 221298 397492
rect 221181 397432 221186 397488
rect 221181 397428 221228 397432
rect 221292 397430 221338 397490
rect 221292 397428 221298 397430
rect 222142 397428 222148 397492
rect 222212 397490 222218 397492
rect 222285 397490 222351 397493
rect 223757 397492 223823 397493
rect 225137 397492 225203 397493
rect 223757 397490 223804 397492
rect 222212 397488 222351 397490
rect 222212 397432 222290 397488
rect 222346 397432 222351 397488
rect 222212 397430 222351 397432
rect 223712 397488 223804 397490
rect 223712 397432 223762 397488
rect 223712 397430 223804 397432
rect 222212 397428 222218 397430
rect 219709 397427 219775 397428
rect 220997 397427 221063 397428
rect 221181 397427 221247 397428
rect 222285 397427 222351 397430
rect 223757 397428 223804 397430
rect 223868 397428 223874 397492
rect 225086 397490 225092 397492
rect 225046 397430 225092 397490
rect 225156 397488 225203 397492
rect 225198 397432 225203 397488
rect 225086 397428 225092 397430
rect 225156 397428 225203 397432
rect 223757 397427 223823 397428
rect 225137 397427 225203 397428
rect 228909 397492 228975 397493
rect 228909 397488 228956 397492
rect 229020 397490 229026 397492
rect 230013 397490 230079 397493
rect 230238 397490 230244 397492
rect 228909 397432 228914 397488
rect 228909 397428 228956 397432
rect 229020 397430 229066 397490
rect 230013 397488 230244 397490
rect 230013 397432 230018 397488
rect 230074 397432 230244 397488
rect 230013 397430 230244 397432
rect 229020 397428 229026 397430
rect 228909 397427 228975 397428
rect 230013 397427 230079 397430
rect 230238 397428 230244 397430
rect 230308 397428 230314 397492
rect 230974 397428 230980 397492
rect 231044 397490 231050 397492
rect 231669 397490 231735 397493
rect 233049 397492 233115 397493
rect 232998 397490 233004 397492
rect 231044 397488 231735 397490
rect 231044 397432 231674 397488
rect 231730 397432 231735 397488
rect 231044 397430 231735 397432
rect 232958 397430 233004 397490
rect 233068 397488 233115 397492
rect 233110 397432 233115 397488
rect 231044 397428 231050 397430
rect 231669 397427 231735 397430
rect 232998 397428 233004 397430
rect 233068 397428 233115 397432
rect 233049 397427 233115 397428
rect 234245 397492 234311 397493
rect 234245 397488 234292 397492
rect 234356 397490 234362 397492
rect 234245 397432 234250 397488
rect 234245 397428 234292 397432
rect 234356 397430 234402 397490
rect 234356 397428 234362 397430
rect 235574 397428 235580 397492
rect 235644 397490 235650 397492
rect 235809 397490 235875 397493
rect 237189 397492 237255 397493
rect 238569 397492 238635 397493
rect 237189 397490 237236 397492
rect 235644 397488 235875 397490
rect 235644 397432 235814 397488
rect 235870 397432 235875 397488
rect 235644 397430 235875 397432
rect 237144 397488 237236 397490
rect 237144 397432 237194 397488
rect 237144 397430 237236 397432
rect 235644 397428 235650 397430
rect 234245 397427 234311 397428
rect 235809 397427 235875 397430
rect 237189 397428 237236 397430
rect 237300 397428 237306 397492
rect 238518 397490 238524 397492
rect 238478 397430 238524 397490
rect 238588 397488 238635 397492
rect 238630 397432 238635 397488
rect 238518 397428 238524 397430
rect 238588 397428 238635 397432
rect 239622 397428 239628 397492
rect 239692 397490 239698 397492
rect 239765 397490 239831 397493
rect 239949 397492 240015 397493
rect 241329 397492 241395 397493
rect 239949 397490 239996 397492
rect 239692 397488 239831 397490
rect 239692 397432 239770 397488
rect 239826 397432 239831 397488
rect 239692 397430 239831 397432
rect 239904 397488 239996 397490
rect 239904 397432 239954 397488
rect 239904 397430 239996 397432
rect 239692 397428 239698 397430
rect 237189 397427 237255 397428
rect 238569 397427 238635 397428
rect 239765 397427 239831 397430
rect 239949 397428 239996 397430
rect 240060 397428 240066 397492
rect 241278 397490 241284 397492
rect 241238 397430 241284 397490
rect 241348 397488 241395 397492
rect 241390 397432 241395 397488
rect 241278 397428 241284 397430
rect 241348 397428 241395 397432
rect 242566 397428 242572 397492
rect 242636 397490 242642 397492
rect 242709 397490 242775 397493
rect 242636 397488 242775 397490
rect 242636 397432 242714 397488
rect 242770 397432 242775 397488
rect 242636 397430 242775 397432
rect 242636 397428 242642 397430
rect 239949 397427 240015 397428
rect 241329 397427 241395 397428
rect 242709 397427 242775 397430
rect 243854 397428 243860 397492
rect 243924 397490 243930 397492
rect 243997 397490 244063 397493
rect 245469 397492 245535 397493
rect 246849 397492 246915 397493
rect 245469 397490 245516 397492
rect 243924 397488 244063 397490
rect 243924 397432 244002 397488
rect 244058 397432 244063 397488
rect 243924 397430 244063 397432
rect 245424 397488 245516 397490
rect 245424 397432 245474 397488
rect 245424 397430 245516 397432
rect 243924 397428 243930 397430
rect 243997 397427 244063 397430
rect 245469 397428 245516 397430
rect 245580 397428 245586 397492
rect 246798 397490 246804 397492
rect 246758 397430 246804 397490
rect 246868 397488 246915 397492
rect 248229 397492 248295 397493
rect 248229 397490 248276 397492
rect 246910 397432 246915 397488
rect 246798 397428 246804 397430
rect 246868 397428 246915 397432
rect 248184 397488 248276 397490
rect 248184 397432 248234 397488
rect 248184 397430 248276 397432
rect 245469 397427 245535 397428
rect 246849 397427 246915 397428
rect 248229 397428 248276 397430
rect 248340 397428 248346 397492
rect 249006 397428 249012 397492
rect 249076 397490 249082 397492
rect 249609 397490 249675 397493
rect 249076 397488 249675 397490
rect 249076 397432 249614 397488
rect 249670 397432 249675 397488
rect 249076 397430 249675 397432
rect 249076 397428 249082 397430
rect 248229 397427 248295 397428
rect 249609 397427 249675 397430
rect 250294 397428 250300 397492
rect 250364 397490 250370 397492
rect 250805 397490 250871 397493
rect 250989 397492 251055 397493
rect 252369 397492 252435 397493
rect 250989 397490 251036 397492
rect 250364 397488 250871 397490
rect 250364 397432 250810 397488
rect 250866 397432 250871 397488
rect 250364 397430 250871 397432
rect 250944 397488 251036 397490
rect 250944 397432 250994 397488
rect 250944 397430 251036 397432
rect 250364 397428 250370 397430
rect 250805 397427 250871 397430
rect 250989 397428 251036 397430
rect 251100 397428 251106 397492
rect 252318 397490 252324 397492
rect 252278 397430 252324 397490
rect 252388 397488 252435 397492
rect 252430 397432 252435 397488
rect 252318 397428 252324 397430
rect 252388 397428 252435 397432
rect 253054 397428 253060 397492
rect 253124 397490 253130 397492
rect 253197 397490 253263 397493
rect 253565 397492 253631 397493
rect 253565 397490 253612 397492
rect 253124 397488 253263 397490
rect 253124 397432 253202 397488
rect 253258 397432 253263 397488
rect 253124 397430 253263 397432
rect 253520 397488 253612 397490
rect 253520 397432 253570 397488
rect 253520 397430 253612 397432
rect 253124 397428 253130 397430
rect 250989 397427 251055 397428
rect 252369 397427 252435 397428
rect 253197 397427 253263 397430
rect 253565 397428 253612 397430
rect 253676 397428 253682 397492
rect 253890 397490 253950 397974
rect 254025 398032 256115 398034
rect 254025 397976 254030 398032
rect 254086 397976 256054 398032
rect 256110 397976 256115 398032
rect 254025 397974 256115 397976
rect 256190 398034 256250 398110
rect 494053 398107 494119 398110
rect 507853 398034 507919 398037
rect 256190 398032 507919 398034
rect 256190 397976 507858 398032
rect 507914 397976 507919 398032
rect 256190 397974 507919 397976
rect 254025 397971 254091 397974
rect 256049 397971 256115 397974
rect 507853 397971 507919 397974
rect 254710 397836 254716 397900
rect 254780 397898 254786 397900
rect 255221 397898 255287 397901
rect 254780 397896 255287 397898
rect 254780 397840 255226 397896
rect 255282 397840 255287 397896
rect 254780 397838 255287 397840
rect 254780 397836 254786 397838
rect 255221 397835 255287 397838
rect 255589 397898 255655 397901
rect 275277 397898 275343 397901
rect 255589 397896 275343 397898
rect 255589 397840 255594 397896
rect 255650 397840 275282 397896
rect 275338 397840 275343 397896
rect 255589 397838 275343 397840
rect 255589 397835 255655 397838
rect 275277 397835 275343 397838
rect 293166 397836 293172 397900
rect 293236 397898 293242 397900
rect 379237 397898 379303 397901
rect 293236 397896 379303 397898
rect 293236 397840 379242 397896
rect 379298 397840 379303 397896
rect 293236 397838 379303 397840
rect 293236 397836 293242 397838
rect 379237 397835 379303 397838
rect 254894 397700 254900 397764
rect 254964 397762 254970 397764
rect 255037 397762 255103 397765
rect 254964 397760 255103 397762
rect 254964 397704 255042 397760
rect 255098 397704 255103 397760
rect 254964 397702 255103 397704
rect 254964 397700 254970 397702
rect 255037 397699 255103 397702
rect 255129 397628 255195 397629
rect 255078 397626 255084 397628
rect 255038 397566 255084 397626
rect 255148 397624 255195 397628
rect 255190 397568 255195 397624
rect 255078 397564 255084 397566
rect 255148 397564 255195 397568
rect 255129 397563 255195 397564
rect 483013 397490 483079 397493
rect 253890 397488 483079 397490
rect 253890 397432 483018 397488
rect 483074 397432 483079 397488
rect 253890 397430 483079 397432
rect 253565 397427 253631 397428
rect 483013 397427 483079 397430
rect 210417 397352 212826 397354
rect 210417 397296 210422 397352
rect 210478 397296 212826 397352
rect 210417 397294 212826 397296
rect 234521 397354 234587 397357
rect 310513 397354 310579 397357
rect 234521 397352 310579 397354
rect 234521 397296 234526 397352
rect 234582 397296 310518 397352
rect 310574 397296 310579 397352
rect 234521 397294 310579 397296
rect 210417 397291 210483 397294
rect 234521 397291 234587 397294
rect 310513 397291 310579 397294
rect 235625 397218 235691 397221
rect 324313 397218 324379 397221
rect 235625 397216 324379 397218
rect 235625 397160 235630 397216
rect 235686 397160 324318 397216
rect 324374 397160 324379 397216
rect 235625 397158 324379 397160
rect 235625 397155 235691 397158
rect 324313 397155 324379 397158
rect 238661 397082 238727 397085
rect 364333 397082 364399 397085
rect 238661 397080 364399 397082
rect 238661 397024 238666 397080
rect 238722 397024 364338 397080
rect 364394 397024 364399 397080
rect 238661 397022 364399 397024
rect 238661 397019 238727 397022
rect 364333 397019 364399 397022
rect 241421 396946 241487 396949
rect 398833 396946 398899 396949
rect 241421 396944 398899 396946
rect 241421 396888 241426 396944
rect 241482 396888 398838 396944
rect 398894 396888 398899 396944
rect 241421 396886 398899 396888
rect 241421 396883 241487 396886
rect 398833 396883 398899 396886
rect 100753 396810 100819 396813
rect 218145 396810 218211 396813
rect 100753 396808 218211 396810
rect 100753 396752 100758 396808
rect 100814 396752 218150 396808
rect 218206 396752 218211 396808
rect 100753 396750 218211 396752
rect 100753 396747 100819 396750
rect 218145 396747 218211 396750
rect 244365 396810 244431 396813
rect 431953 396810 432019 396813
rect 244365 396808 432019 396810
rect 244365 396752 244370 396808
rect 244426 396752 431958 396808
rect 432014 396752 432019 396808
rect 244365 396750 432019 396752
rect 244365 396747 244431 396750
rect 431953 396747 432019 396750
rect 64873 396674 64939 396677
rect 215385 396674 215451 396677
rect 64873 396672 215451 396674
rect 64873 396616 64878 396672
rect 64934 396616 215390 396672
rect 215446 396616 215451 396672
rect 64873 396614 215451 396616
rect 64873 396611 64939 396614
rect 215385 396611 215451 396614
rect 245561 396674 245627 396677
rect 452653 396674 452719 396677
rect 245561 396672 452719 396674
rect 245561 396616 245566 396672
rect 245622 396616 452658 396672
rect 452714 396616 452719 396672
rect 245561 396614 452719 396616
rect 245561 396611 245627 396614
rect 452653 396611 452719 396614
rect 246982 396476 246988 396540
rect 247052 396538 247058 396540
rect 257337 396538 257403 396541
rect 247052 396536 257403 396538
rect 247052 396480 257342 396536
rect 257398 396480 257403 396536
rect 247052 396478 257403 396480
rect 247052 396476 247058 396478
rect 257337 396475 257403 396478
rect 209865 396402 209931 396405
rect 226425 396402 226491 396405
rect 209865 396400 226491 396402
rect 209865 396344 209870 396400
rect 209926 396344 226430 396400
rect 226486 396344 226491 396400
rect 209865 396342 226491 396344
rect 209865 396339 209931 396342
rect 226425 396339 226491 396342
rect 118693 395722 118759 395725
rect 219617 395722 219683 395725
rect 118693 395720 219683 395722
rect 118693 395664 118698 395720
rect 118754 395664 219622 395720
rect 219678 395664 219683 395720
rect 118693 395662 219683 395664
rect 118693 395659 118759 395662
rect 219617 395659 219683 395662
rect 230422 395660 230428 395724
rect 230492 395722 230498 395724
rect 255313 395722 255379 395725
rect 230492 395720 255379 395722
rect 230492 395664 255318 395720
rect 255374 395664 255379 395720
rect 230492 395662 255379 395664
rect 230492 395660 230498 395662
rect 255313 395659 255379 395662
rect 67633 395586 67699 395589
rect 215334 395586 215340 395588
rect 67633 395584 215340 395586
rect 67633 395528 67638 395584
rect 67694 395528 215340 395584
rect 67633 395526 215340 395528
rect 67633 395523 67699 395526
rect 215334 395524 215340 395526
rect 215404 395524 215410 395588
rect 233182 395524 233188 395588
rect 233252 395586 233258 395588
rect 291193 395586 291259 395589
rect 233252 395584 291259 395586
rect 233252 395528 291198 395584
rect 291254 395528 291259 395584
rect 233252 395526 291259 395528
rect 233252 395524 233258 395526
rect 291193 395523 291259 395526
rect 45553 395450 45619 395453
rect 214598 395450 214604 395452
rect 45553 395448 214604 395450
rect 45553 395392 45558 395448
rect 45614 395392 214604 395448
rect 45553 395390 214604 395392
rect 45553 395387 45619 395390
rect 214598 395388 214604 395390
rect 214668 395388 214674 395452
rect 250478 395388 250484 395452
rect 250548 395450 250554 395452
rect 521653 395450 521719 395453
rect 250548 395448 521719 395450
rect 250548 395392 521658 395448
rect 521714 395392 521719 395448
rect 250548 395390 521719 395392
rect 250548 395388 250554 395390
rect 521653 395387 521719 395390
rect 27705 395314 27771 395317
rect 212758 395314 212764 395316
rect 27705 395312 212764 395314
rect 27705 395256 27710 395312
rect 27766 395256 212764 395312
rect 27705 395254 212764 395256
rect 27705 395251 27771 395254
rect 212758 395252 212764 395254
rect 212828 395252 212834 395316
rect 253054 395252 253060 395316
rect 253124 395314 253130 395316
rect 556153 395314 556219 395317
rect 253124 395312 556219 395314
rect 253124 395256 556158 395312
rect 556214 395256 556219 395312
rect 253124 395254 556219 395256
rect 253124 395252 253130 395254
rect 556153 395251 556219 395254
rect 237833 394634 237899 394637
rect 237833 394632 238034 394634
rect 237833 394576 237838 394632
rect 237894 394576 238034 394632
rect 237833 394574 238034 394576
rect 237833 394571 237899 394574
rect 237974 394501 238034 394574
rect 237649 394498 237715 394501
rect 237649 394496 237850 394498
rect 237649 394440 237654 394496
rect 237710 394440 237850 394496
rect 237649 394438 237850 394440
rect 237974 394496 238083 394501
rect 239213 394498 239279 394501
rect 237974 394440 238022 394496
rect 238078 394440 238083 394496
rect 237974 394438 238083 394440
rect 237649 394435 237715 394438
rect 153193 394226 153259 394229
rect 222142 394226 222148 394228
rect 153193 394224 222148 394226
rect 153193 394168 153198 394224
rect 153254 394168 222148 394224
rect 153193 394166 222148 394168
rect 153193 394163 153259 394166
rect 222142 394164 222148 394166
rect 222212 394164 222218 394228
rect 139393 394090 139459 394093
rect 221222 394090 221228 394092
rect 139393 394088 221228 394090
rect 139393 394032 139398 394088
rect 139454 394032 221228 394088
rect 139393 394030 221228 394032
rect 139393 394027 139459 394030
rect 221222 394028 221228 394030
rect 221292 394028 221298 394092
rect 135253 393954 135319 393957
rect 220854 393954 220860 393956
rect 135253 393952 220860 393954
rect 135253 393896 135258 393952
rect 135314 393896 220860 393952
rect 135253 393894 220860 393896
rect 135253 393891 135319 393894
rect 220854 393892 220860 393894
rect 220924 393892 220930 393956
rect 237790 393954 237850 394438
rect 238017 394435 238083 394438
rect 239078 394496 239279 394498
rect 239078 394440 239218 394496
rect 239274 394440 239279 394496
rect 239078 394438 239279 394440
rect 239078 393957 239138 394438
rect 239213 394435 239279 394438
rect 237925 393954 237991 393957
rect 237790 393952 237991 393954
rect 237790 393896 237930 393952
rect 237986 393896 237991 393952
rect 237790 393894 237991 393896
rect 237925 393891 237991 393894
rect 239029 393952 239138 393957
rect 239029 393896 239034 393952
rect 239090 393896 239138 393952
rect 239029 393894 239138 393896
rect 239029 393891 239095 393894
rect 244181 393818 244247 393821
rect 246205 393818 246271 393821
rect 244181 393816 246271 393818
rect 244181 393760 244186 393816
rect 244242 393760 246210 393816
rect 246266 393760 246271 393816
rect 244181 393758 246271 393760
rect 244181 393755 244247 393758
rect 246205 393755 246271 393758
rect 151813 392730 151879 392733
rect 223062 392730 223068 392732
rect 151813 392728 223068 392730
rect 151813 392672 151818 392728
rect 151874 392672 223068 392728
rect 151813 392670 223068 392672
rect 151813 392667 151879 392670
rect 223062 392668 223068 392670
rect 223132 392668 223138 392732
rect 13813 392594 13879 392597
rect 211102 392594 211108 392596
rect 13813 392592 211108 392594
rect 13813 392536 13818 392592
rect 13874 392536 211108 392592
rect 13813 392534 211108 392536
rect 13813 392531 13879 392534
rect 211102 392532 211108 392534
rect 211172 392532 211178 392596
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 253238 355268 253244 355332
rect 253308 355330 253314 355332
rect 557533 355330 557599 355333
rect 253308 355328 557599 355330
rect 253308 355272 557538 355328
rect 557594 355272 557599 355328
rect 253308 355270 557599 355272
rect 253308 355268 253314 355270
rect 557533 355267 557599 355270
rect 230606 354316 230612 354380
rect 230676 354378 230682 354380
rect 273253 354378 273319 354381
rect 230676 354376 273319 354378
rect 230676 354320 273258 354376
rect 273314 354320 273319 354376
rect 230676 354318 273319 354320
rect 230676 354316 230682 354318
rect 273253 354315 273319 354318
rect 247718 354180 247724 354244
rect 247788 354242 247794 354244
rect 488533 354242 488599 354245
rect 247788 354240 488599 354242
rect 247788 354184 488538 354240
rect 488594 354184 488599 354240
rect 247788 354182 488599 354184
rect 247788 354180 247794 354182
rect 488533 354179 488599 354182
rect 102133 354106 102199 354109
rect 218830 354106 218836 354108
rect 102133 354104 218836 354106
rect 102133 354048 102138 354104
rect 102194 354048 218836 354104
rect 102133 354046 218836 354048
rect 102133 354043 102199 354046
rect 218830 354044 218836 354046
rect 218900 354044 218906 354108
rect 251766 354044 251772 354108
rect 251836 354106 251842 354108
rect 538213 354106 538279 354109
rect 251836 354104 538279 354106
rect 251836 354048 538218 354104
rect 538274 354048 538279 354104
rect 251836 354046 538279 354048
rect 251836 354044 251842 354046
rect 538213 354043 538279 354046
rect 84193 353970 84259 353973
rect 217174 353970 217180 353972
rect 84193 353968 217180 353970
rect 84193 353912 84198 353968
rect 84254 353912 217180 353968
rect 84193 353910 217180 353912
rect 84193 353907 84259 353910
rect 217174 353908 217180 353910
rect 217244 353908 217250 353972
rect 253422 353908 253428 353972
rect 253492 353970 253498 353972
rect 558913 353970 558979 353973
rect 253492 353968 558979 353970
rect 253492 353912 558918 353968
rect 558974 353912 558979 353968
rect 253492 353910 558979 353912
rect 253492 353908 253498 353910
rect 558913 353907 558979 353910
rect 238150 352820 238156 352884
rect 238220 352882 238226 352884
rect 360193 352882 360259 352885
rect 238220 352880 360259 352882
rect 238220 352824 360198 352880
rect 360254 352824 360259 352880
rect 238220 352822 360259 352824
rect 238220 352820 238226 352822
rect 360193 352819 360259 352822
rect 248638 352684 248644 352748
rect 248708 352746 248714 352748
rect 506473 352746 506539 352749
rect 248708 352744 506539 352746
rect 248708 352688 506478 352744
rect 506534 352688 506539 352744
rect 248708 352686 506539 352688
rect 248708 352684 248714 352686
rect 506473 352683 506539 352686
rect 191833 352610 191899 352613
rect 225454 352610 225460 352612
rect 191833 352608 225460 352610
rect 191833 352552 191838 352608
rect 191894 352552 225460 352608
rect 191833 352550 225460 352552
rect 191833 352547 191899 352550
rect 225454 352548 225460 352550
rect 225524 352548 225530 352612
rect 254710 352548 254716 352612
rect 254780 352610 254786 352612
rect 576853 352610 576919 352613
rect 254780 352608 576919 352610
rect 254780 352552 576858 352608
rect 576914 352552 576919 352608
rect 254780 352550 576919 352552
rect 254780 352548 254786 352550
rect 576853 352547 576919 352550
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 241278 351052 241284 351116
rect 241348 351114 241354 351116
rect 398925 351114 398991 351117
rect 241348 351112 398991 351114
rect 241348 351056 398930 351112
rect 398986 351056 398991 351112
rect 241348 351054 398991 351056
rect 241348 351052 241354 351054
rect 398925 351051 398991 351054
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect -960 293118 674 293178
rect -960 293042 480 293118
rect 614 293042 674 293118
rect -960 293028 674 293042
rect 246 292982 674 293028
rect 246 292634 306 292982
rect 203374 292634 203380 292636
rect 246 292574 203380 292634
rect 203374 292572 203380 292574
rect 203444 292572 203450 292636
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3969 254146 4035 254149
rect -960 254144 4035 254146
rect -960 254088 3974 254144
rect 4030 254088 4035 254144
rect -960 254086 4035 254088
rect -960 253996 480 254086
rect 3969 254083 4035 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3877 241090 3943 241093
rect -960 241088 3943 241090
rect -960 241032 3882 241088
rect 3938 241032 3943 241088
rect -960 241030 3943 241032
rect -960 240940 480 241030
rect 3877 241027 3943 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3049 214978 3115 214981
rect -960 214976 3115 214978
rect -960 214920 3054 214976
rect 3110 214920 3115 214976
rect -960 214918 3115 214920
rect -960 214828 480 214918
rect 3049 214915 3115 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3785 201922 3851 201925
rect -960 201920 3851 201922
rect -960 201864 3790 201920
rect 3846 201864 3851 201920
rect -960 201862 3851 201864
rect -960 201772 480 201862
rect 3785 201859 3851 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3693 188866 3759 188869
rect -960 188864 3759 188866
rect -960 188808 3698 188864
rect 3754 188808 3759 188864
rect -960 188806 3759 188808
rect -960 188716 480 188806
rect 3693 188803 3759 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 187693 178666 187759 178669
rect 225270 178666 225276 178668
rect 187693 178664 225276 178666
rect 187693 178608 187698 178664
rect 187754 178608 225276 178664
rect 187693 178606 225276 178608
rect 187693 178603 187759 178606
rect 225270 178604 225276 178606
rect 225340 178604 225346 178668
rect 173893 177578 173959 177581
rect 224166 177578 224172 177580
rect 173893 177576 224172 177578
rect 173893 177520 173898 177576
rect 173954 177520 224172 177576
rect 173893 177518 224172 177520
rect 173893 177515 173959 177518
rect 224166 177516 224172 177518
rect 224236 177516 224242 177580
rect 120073 177442 120139 177445
rect 219750 177442 219756 177444
rect 120073 177440 219756 177442
rect 120073 177384 120078 177440
rect 120134 177384 219756 177440
rect 120073 177382 219756 177384
rect 120073 177379 120139 177382
rect 219750 177380 219756 177382
rect 219820 177380 219826 177444
rect 63493 177306 63559 177309
rect 215518 177306 215524 177308
rect 63493 177304 215524 177306
rect 63493 177248 63498 177304
rect 63554 177248 215524 177304
rect 63493 177246 215524 177248
rect 63493 177243 63559 177246
rect 215518 177244 215524 177246
rect 215588 177244 215594 177308
rect 243670 177244 243676 177308
rect 243740 177306 243746 177308
rect 434713 177306 434779 177309
rect 243740 177304 434779 177306
rect 243740 177248 434718 177304
rect 434774 177248 434779 177304
rect 243740 177246 434779 177248
rect 243740 177244 243746 177246
rect 434713 177243 434779 177246
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 251950 86124 251956 86188
rect 252020 86186 252026 86188
rect 539593 86186 539659 86189
rect 252020 86184 539659 86186
rect 252020 86128 539598 86184
rect 539654 86128 539659 86184
rect 252020 86126 539659 86128
rect 252020 86124 252026 86126
rect 539593 86123 539659 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 235206 83404 235212 83468
rect 235276 83466 235282 83468
rect 328453 83466 328519 83469
rect 235276 83464 328519 83466
rect 235276 83408 328458 83464
rect 328514 83408 328519 83464
rect 235276 83406 328519 83408
rect 235276 83404 235282 83406
rect 328453 83403 328519 83406
rect 246430 82044 246436 82108
rect 246500 82106 246506 82108
rect 470593 82106 470659 82109
rect 246500 82104 470659 82106
rect 246500 82048 470598 82104
rect 470654 82048 470659 82104
rect 246500 82046 470659 82048
rect 246500 82044 246506 82046
rect 470593 82043 470659 82046
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 261334 71844 261340 71908
rect 261404 71906 261410 71908
rect 583526 71906 583586 72798
rect 261404 71846 583586 71906
rect 261404 71844 261410 71846
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 190453 46202 190519 46205
rect 225086 46202 225092 46204
rect 190453 46200 225092 46202
rect 190453 46144 190458 46200
rect 190514 46144 225092 46200
rect 190453 46142 225092 46144
rect 190453 46139 190519 46142
rect 225086 46140 225092 46142
rect 225156 46140 225162 46204
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 262438 45596 262444 45660
rect 262508 45658 262514 45660
rect 583526 45658 583586 46142
rect 262508 45598 583586 45658
rect 262508 45596 262514 45598
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 236862 26964 236868 27028
rect 236932 27026 236938 27028
rect 343633 27026 343699 27029
rect 236932 27024 343699 27026
rect 236932 26968 343638 27024
rect 343694 26968 343699 27024
rect 236932 26966 343699 26968
rect 236932 26964 236938 26966
rect 343633 26963 343699 26966
rect 238334 26828 238340 26892
rect 238404 26890 238410 26892
rect 361573 26890 361639 26893
rect 238404 26888 361639 26890
rect 238404 26832 361578 26888
rect 361634 26832 361639 26888
rect 238404 26830 361639 26832
rect 238404 26828 238410 26830
rect 361573 26827 361639 26830
rect 234102 25468 234108 25532
rect 234172 25530 234178 25532
rect 307753 25530 307819 25533
rect 234172 25528 307819 25530
rect 234172 25472 307758 25528
rect 307814 25472 307819 25528
rect 234172 25470 307819 25472
rect 234172 25468 234178 25470
rect 307753 25467 307819 25470
rect 248822 24244 248828 24308
rect 248892 24306 248898 24308
rect 503713 24306 503779 24309
rect 248892 24304 503779 24306
rect 248892 24248 503718 24304
rect 503774 24248 503779 24304
rect 248892 24246 503779 24248
rect 248892 24244 248898 24246
rect 503713 24243 503779 24246
rect 254894 24108 254900 24172
rect 254964 24170 254970 24172
rect 574093 24170 574159 24173
rect 254964 24168 574159 24170
rect 254964 24112 574098 24168
rect 574154 24112 574159 24168
rect 254964 24110 574159 24112
rect 254964 24108 254970 24110
rect 574093 24107 574159 24110
rect 246614 22748 246620 22812
rect 246684 22810 246690 22812
rect 466453 22810 466519 22813
rect 246684 22808 466519 22810
rect 246684 22752 466458 22808
rect 466514 22752 466519 22808
rect 246684 22750 466519 22752
rect 246684 22748 246690 22750
rect 466453 22747 466519 22750
rect 247902 22612 247908 22676
rect 247972 22674 247978 22676
rect 485773 22674 485839 22677
rect 247972 22672 485839 22674
rect 247972 22616 485778 22672
rect 485834 22616 485839 22672
rect 247972 22614 485839 22616
rect 247972 22612 247978 22614
rect 485773 22611 485839 22614
rect 239622 21660 239628 21724
rect 239692 21722 239698 21724
rect 378133 21722 378199 21725
rect 239692 21720 378199 21722
rect 239692 21664 378138 21720
rect 378194 21664 378199 21720
rect 239692 21662 378199 21664
rect 239692 21660 239698 21662
rect 378133 21659 378199 21662
rect 239806 21524 239812 21588
rect 239876 21586 239882 21588
rect 382365 21586 382431 21589
rect 239876 21584 382431 21586
rect 239876 21528 382370 21584
rect 382426 21528 382431 21584
rect 239876 21526 382431 21528
rect 239876 21524 239882 21526
rect 382365 21523 382431 21526
rect 242198 21388 242204 21452
rect 242268 21450 242274 21452
rect 414013 21450 414079 21453
rect 242268 21448 414079 21450
rect 242268 21392 414018 21448
rect 414074 21392 414079 21448
rect 242268 21390 414079 21392
rect 242268 21388 242274 21390
rect 414013 21387 414079 21390
rect 242382 21252 242388 21316
rect 242452 21314 242458 21316
rect 416773 21314 416839 21317
rect 242452 21312 416839 21314
rect 242452 21256 416778 21312
rect 416834 21256 416839 21312
rect 242452 21254 416839 21256
rect 242452 21252 242458 21254
rect 416773 21251 416839 21254
rect 237046 19892 237052 19956
rect 237116 19954 237122 19956
rect 346393 19954 346459 19957
rect 237116 19952 346459 19954
rect 237116 19896 346398 19952
rect 346454 19896 346459 19952
rect 237116 19894 346459 19896
rect 237116 19892 237122 19894
rect 346393 19891 346459 19894
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 295926 19348 295932 19412
rect 295996 19410 296002 19412
rect 583526 19410 583586 19622
rect 295996 19350 583586 19410
rect 295996 19348 296002 19350
rect 232630 18804 232636 18868
rect 232700 18866 232706 18868
rect 289813 18866 289879 18869
rect 232700 18864 289879 18866
rect 232700 18808 289818 18864
rect 289874 18808 289879 18864
rect 232700 18806 289879 18808
rect 232700 18804 232706 18806
rect 289813 18803 289879 18806
rect 232814 18668 232820 18732
rect 232884 18730 232890 18732
rect 292573 18730 292639 18733
rect 232884 18728 292639 18730
rect 232884 18672 292578 18728
rect 292634 18672 292639 18728
rect 232884 18670 292639 18672
rect 232884 18668 232890 18670
rect 292573 18667 292639 18670
rect 234286 18532 234292 18596
rect 234356 18594 234362 18596
rect 307845 18594 307911 18597
rect 234356 18592 307911 18594
rect 234356 18536 307850 18592
rect 307906 18536 307911 18592
rect 234356 18534 307911 18536
rect 234356 18532 234362 18534
rect 307845 18531 307911 18534
rect 243854 16220 243860 16284
rect 243924 16282 243930 16284
rect 432045 16282 432111 16285
rect 243924 16280 432111 16282
rect 243924 16224 432050 16280
rect 432106 16224 432111 16280
rect 243924 16222 432111 16224
rect 243924 16220 243930 16222
rect 432045 16219 432111 16222
rect 250662 16084 250668 16148
rect 250732 16146 250738 16148
rect 523769 16146 523835 16149
rect 250732 16144 523835 16146
rect 250732 16088 523774 16144
rect 523830 16088 523835 16144
rect 250732 16086 523835 16088
rect 250732 16084 250738 16086
rect 523769 16083 523835 16086
rect 170305 16010 170371 16013
rect 223982 16010 223988 16012
rect 170305 16008 223988 16010
rect 170305 15952 170310 16008
rect 170366 15952 223988 16008
rect 170305 15950 223988 15952
rect 170305 15947 170371 15950
rect 223982 15948 223988 15950
rect 224052 15948 224058 16012
rect 252134 15948 252140 16012
rect 252204 16010 252210 16012
rect 541985 16010 542051 16013
rect 252204 16008 542051 16010
rect 252204 15952 541990 16008
rect 542046 15952 542051 16008
rect 252204 15950 542051 15952
rect 252204 15948 252210 15950
rect 541985 15947 542051 15950
rect 99833 15874 99899 15877
rect 218646 15874 218652 15876
rect 99833 15872 218652 15874
rect 99833 15816 99838 15872
rect 99894 15816 218652 15872
rect 99833 15814 218652 15816
rect 99833 15811 99899 15814
rect 218646 15812 218652 15814
rect 218716 15812 218722 15876
rect 253606 15812 253612 15876
rect 253676 15874 253682 15876
rect 556245 15874 556311 15877
rect 253676 15872 556311 15874
rect 253676 15816 556250 15872
rect 556306 15816 556311 15872
rect 253676 15814 556311 15816
rect 253676 15812 253682 15814
rect 556245 15811 556311 15814
rect 138657 14650 138723 14653
rect 216990 14650 216996 14652
rect 138657 14648 216996 14650
rect 138657 14592 138662 14648
rect 138718 14592 216996 14648
rect 138657 14590 216996 14592
rect 138657 14587 138723 14590
rect 216990 14588 216996 14590
rect 217060 14588 217066 14652
rect 50153 14514 50219 14517
rect 214414 14514 214420 14516
rect 50153 14512 214420 14514
rect 50153 14456 50158 14512
rect 50214 14456 214420 14512
rect 50153 14454 214420 14456
rect 50153 14451 50219 14454
rect 214414 14452 214420 14454
rect 214484 14452 214490 14516
rect 250846 14452 250852 14516
rect 250916 14514 250922 14516
rect 520273 14514 520339 14517
rect 250916 14512 520339 14514
rect 250916 14456 520278 14512
rect 520334 14456 520339 14512
rect 250916 14454 520339 14456
rect 250916 14452 250922 14454
rect 520273 14451 520339 14454
rect 88977 13154 89043 13157
rect 211470 13154 211476 13156
rect 88977 13152 211476 13154
rect 88977 13096 88982 13152
rect 89038 13096 211476 13152
rect 88977 13094 211476 13096
rect 88977 13091 89043 13094
rect 211470 13092 211476 13094
rect 211540 13092 211546 13156
rect 246798 13092 246804 13156
rect 246868 13154 246874 13156
rect 469857 13154 469923 13157
rect 246868 13152 469923 13154
rect 246868 13096 469862 13152
rect 469918 13096 469923 13152
rect 246868 13094 469923 13096
rect 246868 13092 246874 13094
rect 469857 13091 469923 13094
rect 66713 13018 66779 13021
rect 215702 13018 215708 13020
rect 66713 13016 215708 13018
rect 66713 12960 66718 13016
rect 66774 12960 215708 13016
rect 66713 12958 215708 12960
rect 66713 12955 66779 12958
rect 215702 12956 215708 12958
rect 215772 12956 215778 13020
rect 248086 12956 248092 13020
rect 248156 13018 248162 13020
rect 484761 13018 484827 13021
rect 248156 13016 484827 13018
rect 248156 12960 484766 13016
rect 484822 12960 484827 13016
rect 248156 12958 484827 12960
rect 248156 12956 248162 12958
rect 484761 12955 484827 12958
rect 122281 12066 122347 12069
rect 219566 12066 219572 12068
rect 122281 12064 219572 12066
rect 122281 12008 122286 12064
rect 122342 12008 219572 12064
rect 122281 12006 219572 12008
rect 122281 12003 122347 12006
rect 219566 12004 219572 12006
rect 219636 12004 219642 12068
rect 48497 11930 48563 11933
rect 214230 11930 214236 11932
rect 48497 11928 214236 11930
rect 48497 11872 48502 11928
rect 48558 11872 214236 11928
rect 48497 11870 214236 11872
rect 48497 11867 48563 11870
rect 214230 11868 214236 11870
rect 214300 11868 214306 11932
rect 30097 11794 30163 11797
rect 212574 11794 212580 11796
rect 30097 11792 212580 11794
rect 30097 11736 30102 11792
rect 30158 11736 212580 11792
rect 30097 11734 212580 11736
rect 30097 11731 30163 11734
rect 212574 11732 212580 11734
rect 212644 11732 212650 11796
rect 244038 11732 244044 11796
rect 244108 11794 244114 11796
rect 433977 11794 434043 11797
rect 244108 11792 434043 11794
rect 244108 11736 433982 11792
rect 434038 11736 434043 11792
rect 244108 11734 434043 11736
rect 244108 11732 244114 11734
rect 433977 11731 434043 11734
rect 17033 11658 17099 11661
rect 211286 11658 211292 11660
rect 17033 11656 211292 11658
rect 17033 11600 17038 11656
rect 17094 11600 211292 11656
rect 17033 11598 211292 11600
rect 17033 11595 17099 11598
rect 211286 11596 211292 11598
rect 211356 11596 211362 11660
rect 245510 11596 245516 11660
rect 245580 11658 245586 11660
rect 451641 11658 451707 11661
rect 245580 11656 451707 11658
rect 245580 11600 451646 11656
rect 451702 11600 451707 11656
rect 245580 11598 451707 11600
rect 245580 11596 245586 11598
rect 451641 11595 451707 11598
rect 185577 10570 185643 10573
rect 219198 10570 219204 10572
rect 185577 10568 219204 10570
rect 185577 10512 185582 10568
rect 185638 10512 219204 10568
rect 185577 10510 219204 10512
rect 185577 10507 185643 10510
rect 219198 10508 219204 10510
rect 219268 10508 219274 10572
rect 239990 10508 239996 10572
rect 240060 10570 240066 10572
rect 381169 10570 381235 10573
rect 240060 10568 381235 10570
rect 240060 10512 381174 10568
rect 381230 10512 381235 10568
rect 240060 10510 381235 10512
rect 240060 10508 240066 10510
rect 381169 10507 381235 10510
rect 86401 10434 86467 10437
rect 216622 10434 216628 10436
rect 86401 10432 216628 10434
rect 86401 10376 86406 10432
rect 86462 10376 216628 10432
rect 86401 10374 216628 10376
rect 86401 10371 86467 10374
rect 216622 10372 216628 10374
rect 216692 10372 216698 10436
rect 242750 10372 242756 10436
rect 242820 10434 242826 10436
rect 412633 10434 412699 10437
rect 242820 10432 412699 10434
rect 242820 10376 412638 10432
rect 412694 10376 412699 10432
rect 242820 10374 412699 10376
rect 242820 10372 242826 10374
rect 412633 10371 412699 10374
rect 83273 10298 83339 10301
rect 216806 10298 216812 10300
rect 83273 10296 216812 10298
rect 83273 10240 83278 10296
rect 83334 10240 216812 10296
rect 83273 10238 216812 10240
rect 83273 10235 83339 10238
rect 216806 10236 216812 10238
rect 216876 10236 216882 10300
rect 242566 10236 242572 10300
rect 242636 10298 242642 10300
rect 415393 10298 415459 10301
rect 242636 10296 415459 10298
rect 242636 10240 415398 10296
rect 415454 10240 415459 10296
rect 242636 10238 415459 10240
rect 242636 10236 242642 10238
rect 415393 10235 415459 10238
rect 88241 9210 88307 9213
rect 211654 9210 211660 9212
rect 88241 9208 211660 9210
rect 88241 9152 88246 9208
rect 88302 9152 211660 9208
rect 88241 9150 211660 9152
rect 88241 9147 88307 9150
rect 211654 9148 211660 9150
rect 211724 9148 211730 9212
rect 1669 9074 1735 9077
rect 209998 9074 210004 9076
rect 1669 9072 210004 9074
rect 1669 9016 1674 9072
rect 1730 9016 210004 9072
rect 1669 9014 210004 9016
rect 1669 9011 1735 9014
rect 209998 9012 210004 9014
rect 210068 9012 210074 9076
rect 235390 9012 235396 9076
rect 235460 9074 235466 9076
rect 326797 9074 326863 9077
rect 235460 9072 326863 9074
rect 235460 9016 326802 9072
rect 326858 9016 326863 9072
rect 235460 9014 326863 9016
rect 235460 9012 235466 9014
rect 326797 9011 326863 9014
rect 565 8938 631 8941
rect 209814 8938 209820 8940
rect 565 8936 209820 8938
rect 565 8880 570 8936
rect 626 8880 209820 8936
rect 565 8878 209820 8880
rect 565 8875 631 8878
rect 209814 8876 209820 8878
rect 209884 8876 209890 8940
rect 238518 8876 238524 8940
rect 238588 8938 238594 8940
rect 363505 8938 363571 8941
rect 238588 8936 363571 8938
rect 238588 8880 363510 8936
rect 363566 8880 363571 8936
rect 238588 8878 363571 8880
rect 238588 8876 238594 8878
rect 363505 8875 363571 8878
rect 138841 7850 138907 7853
rect 221406 7850 221412 7852
rect 138841 7848 221412 7850
rect 138841 7792 138846 7848
rect 138902 7792 221412 7848
rect 138841 7790 221412 7792
rect 138841 7787 138907 7790
rect 221406 7788 221412 7790
rect 221476 7788 221482 7852
rect 137645 7714 137711 7717
rect 221038 7714 221044 7716
rect 137645 7712 221044 7714
rect 137645 7656 137650 7712
rect 137706 7656 221044 7712
rect 137645 7654 221044 7656
rect 137645 7651 137711 7654
rect 221038 7652 221044 7654
rect 221108 7652 221114 7716
rect 233918 7652 233924 7716
rect 233988 7714 233994 7716
rect 310237 7714 310303 7717
rect 233988 7712 310303 7714
rect 233988 7656 310242 7712
rect 310298 7656 310303 7712
rect 233988 7654 310303 7656
rect 233988 7652 233994 7654
rect 310237 7651 310303 7654
rect 51349 7578 51415 7581
rect 214046 7578 214052 7580
rect 51349 7576 214052 7578
rect 51349 7520 51354 7576
rect 51410 7520 214052 7576
rect 51349 7518 214052 7520
rect 51349 7515 51415 7518
rect 214046 7516 214052 7518
rect 214116 7516 214122 7580
rect 235574 7516 235580 7580
rect 235644 7578 235650 7580
rect 327993 7578 328059 7581
rect 235644 7576 328059 7578
rect 235644 7520 327998 7576
rect 328054 7520 328059 7576
rect 235644 7518 328059 7520
rect 235644 7516 235650 7518
rect 327993 7515 328059 7518
rect 230790 6700 230796 6764
rect 230860 6762 230866 6764
rect 276013 6762 276079 6765
rect 230860 6760 276079 6762
rect 230860 6704 276018 6760
rect 276074 6704 276079 6760
rect 230860 6702 276079 6704
rect 230860 6700 230866 6702
rect 276013 6699 276079 6702
rect -960 6490 480 6580
rect 232998 6564 233004 6628
rect 233068 6626 233074 6628
rect 292573 6626 292639 6629
rect 583520 6626 584960 6716
rect 233068 6624 292639 6626
rect 233068 6568 292578 6624
rect 292634 6568 292639 6624
rect 233068 6566 292639 6568
rect 233068 6564 233074 6566
rect 292573 6563 292639 6566
rect 583342 6566 584960 6626
rect 3366 6490 3372 6492
rect -960 6430 3372 6490
rect -960 6340 480 6430
rect 3366 6428 3372 6430
rect 3436 6428 3442 6492
rect 237230 6428 237236 6492
rect 237300 6490 237306 6492
rect 345749 6490 345815 6493
rect 237300 6488 345815 6490
rect 237300 6432 345754 6488
rect 345810 6432 345815 6488
rect 237300 6430 345815 6432
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect 237300 6428 237306 6430
rect 345749 6427 345815 6430
rect 194409 6354 194475 6357
rect 224902 6354 224908 6356
rect 194409 6352 224908 6354
rect 194409 6296 194414 6352
rect 194470 6296 224908 6352
rect 194409 6294 224908 6296
rect 194409 6291 194475 6294
rect 224902 6292 224908 6294
rect 224972 6292 224978 6356
rect 228398 6292 228404 6356
rect 228468 6354 228474 6356
rect 339861 6354 339927 6357
rect 228468 6352 339927 6354
rect 228468 6296 339866 6352
rect 339922 6296 339927 6352
rect 228468 6294 339927 6296
rect 228468 6292 228474 6294
rect 339861 6291 339927 6294
rect 173157 6218 173223 6221
rect 223798 6218 223804 6220
rect 173157 6216 223804 6218
rect 173157 6160 173162 6216
rect 173218 6160 223804 6216
rect 173157 6158 223804 6160
rect 173157 6155 173223 6158
rect 223798 6156 223804 6158
rect 223868 6156 223874 6220
rect 255078 6156 255084 6220
rect 255148 6218 255154 6220
rect 576301 6218 576367 6221
rect 255148 6216 576367 6218
rect 255148 6160 576306 6216
rect 576362 6160 576367 6216
rect 255148 6158 576367 6160
rect 255148 6156 255154 6158
rect 576301 6155 576367 6158
rect 298502 5612 298508 5676
rect 298572 5674 298578 5676
rect 583526 5674 583586 6430
rect 298572 5614 583586 5674
rect 298572 5612 298578 5614
rect 230054 5476 230060 5540
rect 230124 5538 230130 5540
rect 234889 5538 234955 5541
rect 230124 5536 234955 5538
rect 230124 5480 234894 5536
rect 234950 5480 234955 5536
rect 230124 5478 234955 5480
rect 230124 5476 230130 5478
rect 234889 5475 234955 5478
rect 229870 5068 229876 5132
rect 229940 5130 229946 5132
rect 254669 5130 254735 5133
rect 229940 5128 254735 5130
rect 229940 5072 254674 5128
rect 254730 5072 254735 5128
rect 229940 5070 254735 5072
rect 229940 5068 229946 5070
rect 254669 5067 254735 5070
rect 251030 4932 251036 4996
rect 251100 4994 251106 4996
rect 523033 4994 523099 4997
rect 251100 4992 523099 4994
rect 251100 4936 523038 4992
rect 523094 4936 523099 4992
rect 251100 4934 523099 4936
rect 251100 4932 251106 4934
rect 523033 4931 523099 4934
rect 252318 4796 252324 4860
rect 252388 4858 252394 4860
rect 540789 4858 540855 4861
rect 252388 4856 540855 4858
rect 252388 4800 540794 4856
rect 540850 4800 540855 4856
rect 252388 4798 540855 4800
rect 252388 4796 252394 4798
rect 540789 4795 540855 4798
rect 228582 3980 228588 4044
rect 228652 4042 228658 4044
rect 303153 4042 303219 4045
rect 228652 4040 303219 4042
rect 228652 3984 303158 4040
rect 303214 3984 303219 4040
rect 228652 3982 303219 3984
rect 228652 3980 228658 3982
rect 303153 3979 303219 3982
rect 226558 3844 226564 3908
rect 226628 3906 226634 3908
rect 313825 3906 313891 3909
rect 226628 3904 313891 3906
rect 226628 3848 313830 3904
rect 313886 3848 313891 3904
rect 226628 3846 313891 3848
rect 226628 3844 226634 3846
rect 313825 3843 313891 3846
rect 235993 3770 236059 3773
rect 338665 3770 338731 3773
rect 235993 3768 338731 3770
rect 235993 3712 235998 3768
rect 236054 3712 338670 3768
rect 338726 3712 338731 3768
rect 235993 3710 338731 3712
rect 235993 3707 236059 3710
rect 338665 3707 338731 3710
rect 228950 3572 228956 3636
rect 229020 3634 229026 3636
rect 239305 3634 239371 3637
rect 229020 3632 239371 3634
rect 229020 3576 239310 3632
rect 239366 3576 239371 3632
rect 229020 3574 239371 3576
rect 229020 3572 229026 3574
rect 239305 3571 239371 3574
rect 248270 3572 248276 3636
rect 248340 3634 248346 3636
rect 487613 3634 487679 3637
rect 248340 3632 487679 3634
rect 248340 3576 487618 3632
rect 487674 3576 487679 3632
rect 248340 3574 487679 3576
rect 248340 3572 248346 3574
rect 487613 3571 487679 3574
rect 228766 3436 228772 3500
rect 228836 3498 228842 3500
rect 240501 3498 240567 3501
rect 228836 3496 240567 3498
rect 228836 3440 240506 3496
rect 240562 3440 240567 3496
rect 228836 3438 240567 3440
rect 228836 3436 228842 3438
rect 240501 3435 240567 3438
rect 249006 3436 249012 3500
rect 249076 3498 249082 3500
rect 505369 3498 505435 3501
rect 249076 3496 505435 3498
rect 249076 3440 505374 3496
rect 505430 3440 505435 3496
rect 249076 3438 505435 3440
rect 249076 3436 249082 3438
rect 505369 3435 505435 3438
rect 175457 3362 175523 3365
rect 223614 3362 223620 3364
rect 175457 3360 223620 3362
rect 175457 3304 175462 3360
rect 175518 3304 223620 3360
rect 175457 3302 223620 3304
rect 175457 3299 175523 3302
rect 223614 3300 223620 3302
rect 223684 3300 223690 3364
rect 230238 3300 230244 3364
rect 230308 3362 230314 3364
rect 253473 3362 253539 3365
rect 230308 3360 253539 3362
rect 230308 3304 253478 3360
rect 253534 3304 253539 3360
rect 230308 3302 253539 3304
rect 230308 3300 230314 3302
rect 253473 3299 253539 3302
rect 262622 3300 262628 3364
rect 262692 3362 262698 3364
rect 579797 3362 579863 3365
rect 262692 3360 579863 3362
rect 262692 3304 579802 3360
rect 579858 3304 579863 3360
rect 262692 3302 579863 3304
rect 262692 3300 262698 3302
rect 579797 3299 579863 3302
rect 230974 3164 230980 3228
rect 231044 3226 231050 3228
rect 274817 3226 274883 3229
rect 231044 3224 274883 3226
rect 231044 3168 274822 3224
rect 274878 3168 274883 3224
rect 231044 3166 274883 3168
rect 231044 3164 231050 3166
rect 274817 3163 274883 3166
<< via3 >>
rect 102364 597484 102428 597548
rect 110460 597484 110524 597548
rect 207796 597544 207860 597548
rect 207796 597488 207846 597544
rect 207846 597488 207860 597544
rect 207796 597484 207860 597488
rect 208900 597544 208964 597548
rect 208900 597488 208950 597544
rect 208950 597488 208964 597544
rect 208900 597484 208964 597488
rect 210004 597544 210068 597548
rect 210004 597488 210018 597544
rect 210018 597488 210068 597544
rect 210004 597484 210068 597488
rect 211108 597544 211172 597548
rect 211108 597488 211158 597544
rect 211158 597488 211172 597544
rect 211108 597484 211172 597488
rect 212396 597544 212460 597548
rect 212396 597488 212410 597544
rect 212410 597488 212460 597544
rect 212396 597484 212460 597488
rect 213500 597484 213564 597548
rect 214788 597544 214852 597548
rect 214788 597488 214838 597544
rect 214838 597488 214852 597544
rect 214788 597484 214852 597488
rect 215340 597544 215404 597548
rect 215340 597488 215354 597544
rect 215354 597488 215404 597544
rect 215340 597484 215404 597488
rect 215708 597544 215772 597548
rect 215708 597488 215758 597544
rect 215758 597488 215772 597544
rect 215708 597484 215772 597488
rect 225460 597484 225524 597548
rect 235580 597484 235644 597548
rect 245516 597544 245580 597548
rect 245516 597488 245566 597544
rect 245566 597488 245580 597544
rect 245516 597484 245580 597488
rect 250484 597484 250548 597548
rect 317644 597544 317708 597548
rect 317644 597488 317694 597544
rect 317694 597488 317708 597544
rect 317644 597484 317708 597488
rect 320036 597544 320100 597548
rect 320036 597488 320086 597544
rect 320086 597488 320100 597544
rect 320036 597484 320100 597488
rect 321140 597484 321204 597548
rect 322244 597544 322308 597548
rect 322244 597488 322258 597544
rect 322258 597488 322308 597544
rect 322244 597484 322308 597488
rect 323348 597484 323412 597548
rect 325188 597484 325252 597548
rect 325740 597484 325804 597548
rect 330524 597484 330588 597548
rect 345612 597484 345676 597548
rect 360516 597484 360580 597548
rect 440372 597484 440436 597548
rect 450492 597484 450556 597548
rect 460428 597484 460492 597548
rect 92980 597348 93044 597412
rect 99972 597348 100036 597412
rect 318932 597348 318996 597412
rect 324820 597348 324884 597412
rect 335124 597348 335188 597412
rect 428964 597348 429028 597412
rect 430988 597348 431052 597412
rect 435588 597348 435652 597412
rect 98868 597212 98932 597276
rect 104756 597272 104820 597276
rect 104756 597216 104806 597272
rect 104806 597216 104820 597272
rect 104756 597212 104820 597216
rect 230612 597212 230676 597276
rect 314332 597212 314396 597276
rect 422892 597212 422956 597276
rect 427676 597212 427740 597276
rect 94268 597076 94332 597140
rect 101076 597076 101140 597140
rect 205404 597076 205468 597140
rect 350396 597076 350460 597140
rect 433380 597136 433444 597140
rect 433380 597080 433394 597136
rect 433394 597080 433444 597136
rect 433380 597076 433444 597080
rect 434668 597136 434732 597140
rect 434668 597080 434718 597136
rect 434718 597080 434732 597136
rect 434668 597076 434732 597080
rect 103284 596940 103348 597004
rect 105676 596940 105740 597004
rect 130516 596940 130580 597004
rect 340460 596940 340524 597004
rect 424180 596940 424244 597004
rect 429884 596940 429948 597004
rect 431724 596940 431788 597004
rect 97764 596804 97828 596868
rect 105308 596804 105372 596868
rect 240548 596804 240612 596868
rect 315252 596804 315316 596868
rect 465396 596804 465460 596868
rect 125548 596668 125612 596732
rect 435220 596668 435284 596732
rect 445524 596668 445588 596732
rect 135484 596532 135548 596596
rect 140636 596592 140700 596596
rect 140636 596536 140686 596592
rect 140686 596536 140700 596592
rect 140636 596532 140700 596536
rect 312860 596532 312924 596596
rect 202828 596456 202892 596460
rect 202828 596400 202878 596456
rect 202878 596400 202892 596456
rect 202828 596396 202892 596400
rect 425284 596396 425348 596460
rect 95372 596260 95436 596324
rect 115612 596260 115676 596324
rect 120580 596260 120644 596324
rect 204300 596320 204364 596324
rect 204300 596264 204314 596320
rect 204314 596264 204364 596320
rect 204300 596260 204364 596264
rect 219204 596260 219268 596324
rect 354444 596260 354508 596324
rect 455460 596320 455524 596324
rect 455460 596264 455474 596320
rect 455474 596264 455524 596320
rect 455460 596260 455524 596264
rect 470364 596260 470428 596324
rect 282132 589868 282196 589932
rect 407804 526628 407868 526692
rect 408172 523636 408236 523700
rect 408172 489772 408236 489836
rect 92980 488472 93044 488476
rect 92980 488416 92994 488472
rect 92994 488416 93044 488472
rect 92980 488412 93044 488416
rect 94268 488472 94332 488476
rect 94268 488416 94282 488472
rect 94282 488416 94332 488472
rect 94268 488412 94332 488416
rect 95372 488472 95436 488476
rect 95372 488416 95386 488472
rect 95386 488416 95436 488472
rect 95372 488412 95436 488416
rect 97764 488472 97828 488476
rect 97764 488416 97814 488472
rect 97814 488416 97828 488472
rect 97764 488412 97828 488416
rect 98868 488472 98932 488476
rect 98868 488416 98918 488472
rect 98918 488416 98932 488472
rect 98868 488412 98932 488416
rect 99972 488472 100036 488476
rect 99972 488416 100022 488472
rect 100022 488416 100036 488472
rect 99972 488412 100036 488416
rect 101076 488472 101140 488476
rect 101076 488416 101126 488472
rect 101126 488416 101140 488472
rect 101076 488412 101140 488416
rect 102364 488472 102428 488476
rect 102364 488416 102414 488472
rect 102414 488416 102428 488472
rect 102364 488412 102428 488416
rect 104756 488472 104820 488476
rect 104756 488416 104806 488472
rect 104806 488416 104820 488472
rect 104756 488412 104820 488416
rect 105676 488472 105740 488476
rect 105676 488416 105726 488472
rect 105726 488416 105740 488472
rect 105676 488412 105740 488416
rect 204300 488412 204364 488476
rect 214788 488472 214852 488476
rect 214788 488416 214838 488472
rect 214838 488416 214852 488472
rect 214788 488412 214852 488416
rect 211108 488336 211172 488340
rect 211108 488280 211158 488336
rect 211158 488280 211172 488336
rect 211108 488276 211172 488280
rect 213500 488276 213564 488340
rect 215708 488336 215772 488340
rect 215708 488280 215758 488336
rect 215758 488280 215772 488336
rect 215708 488276 215772 488280
rect 314332 488472 314396 488476
rect 314332 488416 314346 488472
rect 314346 488416 314396 488472
rect 314332 488412 314396 488416
rect 315436 488472 315500 488476
rect 315436 488416 315450 488472
rect 315450 488416 315500 488472
rect 315436 488412 315500 488416
rect 422892 488412 422956 488476
rect 424180 488412 424244 488476
rect 425284 488412 425348 488476
rect 105308 488140 105372 488204
rect 110460 488140 110524 488204
rect 203012 488140 203076 488204
rect 465396 488276 465460 488340
rect 429884 488140 429948 488204
rect 435588 488140 435652 488204
rect 407804 488004 407868 488068
rect 103284 487868 103348 487932
rect 208900 487928 208964 487932
rect 208900 487872 208914 487928
rect 208914 487872 208964 487928
rect 208900 487868 208964 487872
rect 313044 487928 313108 487932
rect 313044 487872 313058 487928
rect 313058 487872 313108 487928
rect 313044 487868 313108 487872
rect 324636 487868 324700 487932
rect 325740 487732 325804 487796
rect 430988 487732 431052 487796
rect 427676 487596 427740 487660
rect 428964 487596 429028 487660
rect 212212 487460 212276 487524
rect 320036 487520 320100 487524
rect 320036 487464 320050 487520
rect 320050 487464 320100 487520
rect 320036 487460 320100 487464
rect 323348 487460 323412 487524
rect 433380 487520 433444 487524
rect 433380 487464 433394 487520
rect 433394 487464 433444 487520
rect 433380 487460 433444 487464
rect 322244 487384 322308 487388
rect 322244 487328 322258 487384
rect 322258 487328 322308 487384
rect 322244 487324 322308 487328
rect 432276 487324 432340 487388
rect 434852 487324 434916 487388
rect 115612 487188 115676 487252
rect 120580 487188 120644 487252
rect 125548 487188 125612 487252
rect 130516 487188 130580 487252
rect 135484 487188 135548 487252
rect 140636 487248 140700 487252
rect 140636 487192 140686 487248
rect 140686 487192 140700 487248
rect 140636 487188 140700 487192
rect 203012 487188 203076 487252
rect 205404 487188 205468 487252
rect 207612 487248 207676 487252
rect 207612 487192 207662 487248
rect 207662 487192 207676 487248
rect 207612 487188 207676 487192
rect 210004 487188 210068 487252
rect 215340 487188 215404 487252
rect 220492 487188 220556 487252
rect 225460 487188 225524 487252
rect 230612 487188 230676 487252
rect 235580 487188 235644 487252
rect 240548 487188 240612 487252
rect 245516 487188 245580 487252
rect 250484 487188 250548 487252
rect 317644 487188 317708 487252
rect 318932 487188 318996 487252
rect 321140 487188 321204 487252
rect 325188 487188 325252 487252
rect 330524 487188 330588 487252
rect 335492 487188 335556 487252
rect 340460 487188 340524 487252
rect 345612 487188 345676 487252
rect 350396 487188 350460 487252
rect 355548 487188 355612 487252
rect 360516 487188 360580 487252
rect 435220 487188 435284 487252
rect 440372 487188 440436 487252
rect 445524 487188 445588 487252
rect 450492 487188 450556 487252
rect 455460 487248 455524 487252
rect 455460 487192 455474 487248
rect 455474 487192 455524 487248
rect 455460 487188 455524 487192
rect 460428 487188 460492 487252
rect 470732 487188 470796 487252
rect 382228 454276 382292 454340
rect 382412 454140 382476 454204
rect 293172 448700 293236 448764
rect 3372 446660 3436 446724
rect 258580 446524 258644 446588
rect 282132 446388 282196 446452
rect 298508 446116 298572 446180
rect 264100 445844 264164 445908
rect 262628 445708 262692 445772
rect 262444 444756 262508 444820
rect 261524 444348 261588 444412
rect 260052 444212 260116 444276
rect 209636 444076 209700 444140
rect 210740 444076 210804 444140
rect 238156 444076 238220 444140
rect 256372 444136 256436 444140
rect 256372 444080 256422 444136
rect 256422 444080 256436 444136
rect 256372 444076 256436 444080
rect 245516 444000 245580 444004
rect 245516 443944 245530 444000
rect 245530 443944 245580 444000
rect 245516 443940 245580 443944
rect 251036 444000 251100 444004
rect 251036 443944 251050 444000
rect 251050 443944 251100 444000
rect 251036 443940 251100 443944
rect 220124 443668 220188 443732
rect 261340 443532 261404 443596
rect 203380 442988 203444 443052
rect 220124 442988 220188 443052
rect 251036 442716 251100 442780
rect 245516 442580 245580 442644
rect 238156 442444 238220 442508
rect 210740 442308 210804 442372
rect 209636 442172 209700 442236
rect 295932 442172 295996 442236
rect 256372 441628 256436 441692
rect 260236 441628 260300 441692
rect 383332 425716 383396 425780
rect 383332 412524 383396 412588
rect 383332 402868 383396 402932
rect 260052 401508 260116 401572
rect 383332 401508 383396 401572
rect 252876 399876 252940 399940
rect 214604 398652 214668 398716
rect 205588 398380 205652 398444
rect 211292 398244 211356 398308
rect 205588 398108 205652 398172
rect 252692 399196 252756 399260
rect 250300 398788 250364 398852
rect 252692 398848 252756 398852
rect 252692 398792 252706 398848
rect 252706 398792 252756 398848
rect 252692 398788 252756 398792
rect 252876 398652 252940 398716
rect 258580 398924 258644 398988
rect 264100 398788 264164 398852
rect 228588 398516 228652 398580
rect 253428 398380 253492 398444
rect 246988 398244 247052 398308
rect 216628 397836 216692 397900
rect 223988 397836 224052 397900
rect 224908 397836 224972 397900
rect 228772 397836 228836 397900
rect 211660 397700 211724 397764
rect 212764 397700 212828 397764
rect 214052 397700 214116 397764
rect 215340 397700 215404 397764
rect 216996 397700 217060 397764
rect 223068 397700 223132 397764
rect 224172 397700 224236 397764
rect 225276 397700 225340 397764
rect 228404 397700 228468 397764
rect 260236 398652 260300 398716
rect 261524 398516 261588 398580
rect 230428 397972 230492 398036
rect 233188 397972 233252 398036
rect 209820 397564 209884 397628
rect 211292 397564 211356 397628
rect 210004 397428 210068 397492
rect 211476 397428 211540 397492
rect 212580 397488 212644 397492
rect 214420 397564 214484 397628
rect 215708 397564 215772 397628
rect 217180 397564 217244 397628
rect 218836 397564 218900 397628
rect 219572 397564 219636 397628
rect 220860 397624 220924 397628
rect 220860 397568 220910 397624
rect 220910 397568 220924 397624
rect 220860 397564 220924 397568
rect 221412 397564 221476 397628
rect 223620 397564 223684 397628
rect 225460 397564 225524 397628
rect 226564 397564 226628 397628
rect 242388 397836 242452 397900
rect 247724 397836 247788 397900
rect 250484 397836 250548 397900
rect 251772 397836 251836 397900
rect 230060 397700 230124 397764
rect 230612 397700 230676 397764
rect 232820 397700 232884 397764
rect 233924 397700 233988 397764
rect 235212 397700 235276 397764
rect 236868 397700 236932 397764
rect 238156 397700 238220 397764
rect 242204 397700 242268 397764
rect 243676 397700 243740 397764
rect 246436 397700 246500 397764
rect 247908 397700 247972 397764
rect 248644 397700 248708 397764
rect 250668 397700 250732 397764
rect 251956 397700 252020 397764
rect 253244 397700 253308 397764
rect 229876 397564 229940 397628
rect 230796 397564 230860 397628
rect 232636 397564 232700 397628
rect 234108 397564 234172 397628
rect 235396 397564 235460 397628
rect 237052 397564 237116 397628
rect 238340 397564 238404 397628
rect 239812 397564 239876 397628
rect 242756 397564 242820 397628
rect 244044 397624 244108 397628
rect 244044 397568 244094 397624
rect 244094 397568 244108 397624
rect 244044 397564 244108 397568
rect 246620 397624 246684 397628
rect 246620 397568 246670 397624
rect 246670 397568 246684 397624
rect 246620 397564 246684 397568
rect 248092 397624 248156 397628
rect 248092 397568 248106 397624
rect 248106 397568 248156 397624
rect 248092 397564 248156 397568
rect 248828 397564 248892 397628
rect 250852 397624 250916 397628
rect 250852 397568 250866 397624
rect 250866 397568 250916 397624
rect 250852 397564 250916 397568
rect 252140 397564 252204 397628
rect 212580 397432 212630 397488
rect 212630 397432 212644 397488
rect 212580 397428 212644 397432
rect 214236 397428 214300 397492
rect 215524 397428 215588 397492
rect 216812 397488 216876 397492
rect 216812 397432 216826 397488
rect 216826 397432 216876 397488
rect 216812 397428 216876 397432
rect 218652 397428 218716 397492
rect 219388 397428 219452 397492
rect 219756 397488 219820 397492
rect 219756 397432 219770 397488
rect 219770 397432 219820 397488
rect 219756 397428 219820 397432
rect 221044 397488 221108 397492
rect 221044 397432 221058 397488
rect 221058 397432 221108 397488
rect 221044 397428 221108 397432
rect 221228 397488 221292 397492
rect 221228 397432 221242 397488
rect 221242 397432 221292 397488
rect 221228 397428 221292 397432
rect 222148 397428 222212 397492
rect 223804 397488 223868 397492
rect 223804 397432 223818 397488
rect 223818 397432 223868 397488
rect 223804 397428 223868 397432
rect 225092 397488 225156 397492
rect 225092 397432 225142 397488
rect 225142 397432 225156 397488
rect 225092 397428 225156 397432
rect 228956 397488 229020 397492
rect 228956 397432 228970 397488
rect 228970 397432 229020 397488
rect 228956 397428 229020 397432
rect 230244 397428 230308 397492
rect 230980 397428 231044 397492
rect 233004 397488 233068 397492
rect 233004 397432 233054 397488
rect 233054 397432 233068 397488
rect 233004 397428 233068 397432
rect 234292 397488 234356 397492
rect 234292 397432 234306 397488
rect 234306 397432 234356 397488
rect 234292 397428 234356 397432
rect 235580 397428 235644 397492
rect 237236 397488 237300 397492
rect 237236 397432 237250 397488
rect 237250 397432 237300 397488
rect 237236 397428 237300 397432
rect 238524 397488 238588 397492
rect 238524 397432 238574 397488
rect 238574 397432 238588 397488
rect 238524 397428 238588 397432
rect 239628 397428 239692 397492
rect 239996 397488 240060 397492
rect 239996 397432 240010 397488
rect 240010 397432 240060 397488
rect 239996 397428 240060 397432
rect 241284 397488 241348 397492
rect 241284 397432 241334 397488
rect 241334 397432 241348 397488
rect 241284 397428 241348 397432
rect 242572 397428 242636 397492
rect 243860 397428 243924 397492
rect 245516 397488 245580 397492
rect 245516 397432 245530 397488
rect 245530 397432 245580 397488
rect 245516 397428 245580 397432
rect 246804 397488 246868 397492
rect 246804 397432 246854 397488
rect 246854 397432 246868 397488
rect 246804 397428 246868 397432
rect 248276 397488 248340 397492
rect 248276 397432 248290 397488
rect 248290 397432 248340 397488
rect 248276 397428 248340 397432
rect 249012 397428 249076 397492
rect 250300 397428 250364 397492
rect 251036 397488 251100 397492
rect 251036 397432 251050 397488
rect 251050 397432 251100 397488
rect 251036 397428 251100 397432
rect 252324 397488 252388 397492
rect 252324 397432 252374 397488
rect 252374 397432 252388 397488
rect 252324 397428 252388 397432
rect 253060 397428 253124 397492
rect 253612 397488 253676 397492
rect 253612 397432 253626 397488
rect 253626 397432 253676 397488
rect 253612 397428 253676 397432
rect 254716 397836 254780 397900
rect 293172 397836 293236 397900
rect 254900 397700 254964 397764
rect 255084 397624 255148 397628
rect 255084 397568 255134 397624
rect 255134 397568 255148 397624
rect 255084 397564 255148 397568
rect 246988 396476 247052 396540
rect 230428 395660 230492 395724
rect 215340 395524 215404 395588
rect 233188 395524 233252 395588
rect 214604 395388 214668 395452
rect 250484 395388 250548 395452
rect 212764 395252 212828 395316
rect 253060 395252 253124 395316
rect 222148 394164 222212 394228
rect 221228 394028 221292 394092
rect 220860 393892 220924 393956
rect 223068 392668 223132 392732
rect 211108 392532 211172 392596
rect 253244 355268 253308 355332
rect 230612 354316 230676 354380
rect 247724 354180 247788 354244
rect 218836 354044 218900 354108
rect 251772 354044 251836 354108
rect 217180 353908 217244 353972
rect 253428 353908 253492 353972
rect 238156 352820 238220 352884
rect 248644 352684 248708 352748
rect 225460 352548 225524 352612
rect 254716 352548 254780 352612
rect 241284 351052 241348 351116
rect 203380 292572 203444 292636
rect 225276 178604 225340 178668
rect 224172 177516 224236 177580
rect 219756 177380 219820 177444
rect 215524 177244 215588 177308
rect 243676 177244 243740 177308
rect 251956 86124 252020 86188
rect 235212 83404 235276 83468
rect 246436 82044 246500 82108
rect 261340 71844 261404 71908
rect 225092 46140 225156 46204
rect 262444 45596 262508 45660
rect 236868 26964 236932 27028
rect 238340 26828 238404 26892
rect 234108 25468 234172 25532
rect 248828 24244 248892 24308
rect 254900 24108 254964 24172
rect 246620 22748 246684 22812
rect 247908 22612 247972 22676
rect 239628 21660 239692 21724
rect 239812 21524 239876 21588
rect 242204 21388 242268 21452
rect 242388 21252 242452 21316
rect 237052 19892 237116 19956
rect 295932 19348 295996 19412
rect 232636 18804 232700 18868
rect 232820 18668 232884 18732
rect 234292 18532 234356 18596
rect 243860 16220 243924 16284
rect 250668 16084 250732 16148
rect 223988 15948 224052 16012
rect 252140 15948 252204 16012
rect 218652 15812 218716 15876
rect 253612 15812 253676 15876
rect 216996 14588 217060 14652
rect 214420 14452 214484 14516
rect 250852 14452 250916 14516
rect 211476 13092 211540 13156
rect 246804 13092 246868 13156
rect 215708 12956 215772 13020
rect 248092 12956 248156 13020
rect 219572 12004 219636 12068
rect 214236 11868 214300 11932
rect 212580 11732 212644 11796
rect 244044 11732 244108 11796
rect 211292 11596 211356 11660
rect 245516 11596 245580 11660
rect 219204 10508 219268 10572
rect 239996 10508 240060 10572
rect 216628 10372 216692 10436
rect 242756 10372 242820 10436
rect 216812 10236 216876 10300
rect 242572 10236 242636 10300
rect 211660 9148 211724 9212
rect 210004 9012 210068 9076
rect 235396 9012 235460 9076
rect 209820 8876 209884 8940
rect 238524 8876 238588 8940
rect 221412 7788 221476 7852
rect 221044 7652 221108 7716
rect 233924 7652 233988 7716
rect 214052 7516 214116 7580
rect 235580 7516 235644 7580
rect 230796 6700 230860 6764
rect 233004 6564 233068 6628
rect 3372 6428 3436 6492
rect 237236 6428 237300 6492
rect 224908 6292 224972 6356
rect 228404 6292 228468 6356
rect 223804 6156 223868 6220
rect 255084 6156 255148 6220
rect 298508 5612 298572 5676
rect 230060 5476 230124 5540
rect 229876 5068 229940 5132
rect 251036 4932 251100 4996
rect 252324 4796 252388 4860
rect 228588 3980 228652 4044
rect 226564 3844 226628 3908
rect 228956 3572 229020 3636
rect 248276 3572 248340 3636
rect 228772 3436 228836 3500
rect 249012 3436 249076 3500
rect 223620 3300 223684 3364
rect 230244 3300 230308 3364
rect 262628 3300 262692 3364
rect 230980 3164 231044 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 3371 446724 3437 446725
rect 3371 446660 3372 446724
rect 3436 446660 3437 446724
rect 3371 446659 3437 446660
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 6493 3434 446659
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 3371 6492 3437 6493
rect 3371 6428 3372 6492
rect 3436 6428 3437 6492
rect 3371 6427 3437 6428
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 691292 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 691292 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 691292 87914 700398
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 691292 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 691292 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 691292 123914 700398
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 691292 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 691292 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 691292 159914 700398
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 80952 687454 81300 687486
rect 80952 687218 81008 687454
rect 81244 687218 81300 687454
rect 80952 687134 81300 687218
rect 80952 686898 81008 687134
rect 81244 686898 81300 687134
rect 80952 686866 81300 686898
rect 169760 687454 170108 687486
rect 169760 687218 169816 687454
rect 170052 687218 170108 687454
rect 169760 687134 170108 687218
rect 169760 686898 169816 687134
rect 170052 686898 170108 687134
rect 169760 686866 170108 686898
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 80272 655954 80620 655986
rect 80272 655718 80328 655954
rect 80564 655718 80620 655954
rect 80272 655634 80620 655718
rect 80272 655398 80328 655634
rect 80564 655398 80620 655634
rect 80272 655366 80620 655398
rect 170440 655954 170788 655986
rect 170440 655718 170496 655954
rect 170732 655718 170788 655954
rect 170440 655634 170788 655718
rect 170440 655398 170496 655634
rect 170732 655398 170788 655634
rect 170440 655366 170788 655398
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 80952 651454 81300 651486
rect 80952 651218 81008 651454
rect 81244 651218 81300 651454
rect 80952 651134 81300 651218
rect 80952 650898 81008 651134
rect 81244 650898 81300 651134
rect 80952 650866 81300 650898
rect 169760 651454 170108 651486
rect 169760 651218 169816 651454
rect 170052 651218 170108 651454
rect 169760 651134 170108 651218
rect 169760 650898 169816 651134
rect 170052 650898 170108 651134
rect 169760 650866 170108 650898
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 80272 619954 80620 619986
rect 80272 619718 80328 619954
rect 80564 619718 80620 619954
rect 80272 619634 80620 619718
rect 80272 619398 80328 619634
rect 80564 619398 80620 619634
rect 80272 619366 80620 619398
rect 170440 619954 170788 619986
rect 170440 619718 170496 619954
rect 170732 619718 170788 619954
rect 170440 619634 170788 619718
rect 170440 619398 170496 619634
rect 170732 619398 170788 619634
rect 170440 619366 170788 619398
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 80952 615454 81300 615486
rect 80952 615218 81008 615454
rect 81244 615218 81300 615454
rect 80952 615134 81300 615218
rect 80952 614898 81008 615134
rect 81244 614898 81300 615134
rect 80952 614866 81300 614898
rect 169760 615454 170108 615486
rect 169760 615218 169816 615454
rect 170052 615218 170108 615454
rect 169760 615134 170108 615218
rect 169760 614898 169816 615134
rect 170052 614898 170108 615134
rect 169760 614866 170108 614898
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 92928 599450 92988 600100
rect 94288 599450 94348 600100
rect 95376 599450 95436 600100
rect 92928 599390 93042 599450
rect 92982 597413 93042 599390
rect 94270 599390 94348 599450
rect 95374 599390 95436 599450
rect 97688 599450 97748 600100
rect 98912 599450 98972 600100
rect 100000 599450 100060 600100
rect 101088 599450 101148 600100
rect 97688 599390 97826 599450
rect 92979 597412 93045 597413
rect 92979 597348 92980 597412
rect 93044 597348 93045 597412
rect 92979 597347 93045 597348
rect 94270 597141 94330 599390
rect 94267 597140 94333 597141
rect 94267 597076 94268 597140
rect 94332 597076 94333 597140
rect 94267 597075 94333 597076
rect 95374 596325 95434 599390
rect 97766 596869 97826 599390
rect 98870 599390 98972 599450
rect 99974 599390 100060 599450
rect 101078 599390 101148 599450
rect 102312 599450 102372 600100
rect 103400 599450 103460 600100
rect 104760 599450 104820 600100
rect 102312 599390 102426 599450
rect 98870 597277 98930 599390
rect 99974 597413 100034 599390
rect 99971 597412 100037 597413
rect 99971 597348 99972 597412
rect 100036 597348 100037 597412
rect 99971 597347 100037 597348
rect 98867 597276 98933 597277
rect 98867 597212 98868 597276
rect 98932 597212 98933 597276
rect 98867 597211 98933 597212
rect 101078 597141 101138 599390
rect 102366 597549 102426 599390
rect 103286 599390 103460 599450
rect 104758 599390 104820 599450
rect 105304 599450 105364 600100
rect 105712 599450 105772 600100
rect 110472 599450 110532 600100
rect 105304 599390 105370 599450
rect 102363 597548 102429 597549
rect 102363 597484 102364 597548
rect 102428 597484 102429 597548
rect 102363 597483 102429 597484
rect 101075 597140 101141 597141
rect 101075 597076 101076 597140
rect 101140 597076 101141 597140
rect 101075 597075 101141 597076
rect 103286 597005 103346 599390
rect 104758 597277 104818 599390
rect 104755 597276 104821 597277
rect 104755 597212 104756 597276
rect 104820 597212 104821 597276
rect 104755 597211 104821 597212
rect 103283 597004 103349 597005
rect 103283 596940 103284 597004
rect 103348 596940 103349 597004
rect 103283 596939 103349 596940
rect 105310 596869 105370 599390
rect 105678 599390 105772 599450
rect 110462 599390 110532 599450
rect 115504 599450 115564 600100
rect 120536 599450 120596 600100
rect 125568 599450 125628 600100
rect 115504 599390 115674 599450
rect 120536 599390 120642 599450
rect 105678 597005 105738 599390
rect 110462 597549 110522 599390
rect 110459 597548 110525 597549
rect 110459 597484 110460 597548
rect 110524 597484 110525 597548
rect 110459 597483 110525 597484
rect 105675 597004 105741 597005
rect 105675 596940 105676 597004
rect 105740 596940 105741 597004
rect 105675 596939 105741 596940
rect 97763 596868 97829 596869
rect 97763 596804 97764 596868
rect 97828 596804 97829 596868
rect 97763 596803 97829 596804
rect 105307 596868 105373 596869
rect 105307 596804 105308 596868
rect 105372 596804 105373 596868
rect 105307 596803 105373 596804
rect 115614 596325 115674 599390
rect 120582 596325 120642 599390
rect 125550 599390 125628 599450
rect 130464 599450 130524 600100
rect 135496 599450 135556 600100
rect 130464 599390 130578 599450
rect 125550 596733 125610 599390
rect 130518 597005 130578 599390
rect 135486 599390 135556 599450
rect 140528 599450 140588 600100
rect 140528 599390 140698 599450
rect 130515 597004 130581 597005
rect 130515 596940 130516 597004
rect 130580 596940 130581 597004
rect 130515 596939 130581 596940
rect 125547 596732 125613 596733
rect 125547 596668 125548 596732
rect 125612 596668 125613 596732
rect 125547 596667 125613 596668
rect 135486 596597 135546 599390
rect 140638 596597 140698 599390
rect 135483 596596 135549 596597
rect 135483 596532 135484 596596
rect 135548 596532 135549 596596
rect 135483 596531 135549 596532
rect 140635 596596 140701 596597
rect 140635 596532 140636 596596
rect 140700 596532 140701 596596
rect 140635 596531 140701 596532
rect 95371 596324 95437 596325
rect 95371 596260 95372 596324
rect 95436 596260 95437 596324
rect 95371 596259 95437 596260
rect 115611 596324 115677 596325
rect 115611 596260 115612 596324
rect 115676 596260 115677 596324
rect 115611 596259 115677 596260
rect 120579 596324 120645 596325
rect 120579 596260 120580 596324
rect 120644 596260 120645 596324
rect 120579 596259 120645 596260
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 80272 547954 80620 547986
rect 80272 547718 80328 547954
rect 80564 547718 80620 547954
rect 80272 547634 80620 547718
rect 80272 547398 80328 547634
rect 80564 547398 80620 547634
rect 80272 547366 80620 547398
rect 170440 547954 170788 547986
rect 170440 547718 170496 547954
rect 170732 547718 170788 547954
rect 170440 547634 170788 547718
rect 170440 547398 170496 547634
rect 170732 547398 170788 547634
rect 170440 547366 170788 547398
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 80952 543454 81300 543486
rect 80952 543218 81008 543454
rect 81244 543218 81300 543454
rect 80952 543134 81300 543218
rect 80952 542898 81008 543134
rect 81244 542898 81300 543134
rect 80952 542866 81300 542898
rect 169760 543454 170108 543486
rect 169760 543218 169816 543454
rect 170052 543218 170108 543454
rect 169760 543134 170108 543218
rect 169760 542898 169816 543134
rect 170052 542898 170108 543134
rect 169760 542866 170108 542898
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 80272 511954 80620 511986
rect 80272 511718 80328 511954
rect 80564 511718 80620 511954
rect 80272 511634 80620 511718
rect 80272 511398 80328 511634
rect 80564 511398 80620 511634
rect 80272 511366 80620 511398
rect 170440 511954 170788 511986
rect 170440 511718 170496 511954
rect 170732 511718 170788 511954
rect 170440 511634 170788 511718
rect 170440 511398 170496 511634
rect 170732 511398 170788 511634
rect 170440 511366 170788 511398
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 80952 507454 81300 507486
rect 80952 507218 81008 507454
rect 81244 507218 81300 507454
rect 80952 507134 81300 507218
rect 80952 506898 81008 507134
rect 81244 506898 81300 507134
rect 80952 506866 81300 506898
rect 169760 507454 170108 507486
rect 169760 507218 169816 507454
rect 170052 507218 170108 507454
rect 169760 507134 170108 507218
rect 169760 506898 169816 507134
rect 170052 506898 170108 507134
rect 169760 506866 170108 506898
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 92928 489930 92988 490106
rect 94288 489930 94348 490106
rect 95376 489930 95436 490106
rect 92928 489870 93042 489930
rect 92982 488477 93042 489870
rect 94270 489870 94348 489930
rect 95374 489870 95436 489930
rect 97688 489930 97748 490106
rect 98912 489930 98972 490106
rect 100000 489930 100060 490106
rect 101088 489930 101148 490106
rect 97688 489870 97826 489930
rect 94270 488477 94330 489870
rect 95374 488477 95434 489870
rect 97766 488477 97826 489870
rect 98870 489870 98972 489930
rect 99974 489870 100060 489930
rect 101078 489870 101148 489930
rect 102312 489930 102372 490106
rect 103400 489930 103460 490106
rect 104760 489930 104820 490106
rect 102312 489870 102426 489930
rect 98870 488477 98930 489870
rect 99974 488477 100034 489870
rect 101078 488477 101138 489870
rect 102366 488477 102426 489870
rect 103286 489870 103460 489930
rect 104758 489870 104820 489930
rect 105304 489930 105364 490106
rect 105712 489930 105772 490106
rect 110472 489930 110532 490106
rect 105304 489870 105370 489930
rect 92979 488476 93045 488477
rect 92979 488412 92980 488476
rect 93044 488412 93045 488476
rect 92979 488411 93045 488412
rect 94267 488476 94333 488477
rect 94267 488412 94268 488476
rect 94332 488412 94333 488476
rect 94267 488411 94333 488412
rect 95371 488476 95437 488477
rect 95371 488412 95372 488476
rect 95436 488412 95437 488476
rect 95371 488411 95437 488412
rect 97763 488476 97829 488477
rect 97763 488412 97764 488476
rect 97828 488412 97829 488476
rect 97763 488411 97829 488412
rect 98867 488476 98933 488477
rect 98867 488412 98868 488476
rect 98932 488412 98933 488476
rect 98867 488411 98933 488412
rect 99971 488476 100037 488477
rect 99971 488412 99972 488476
rect 100036 488412 100037 488476
rect 99971 488411 100037 488412
rect 101075 488476 101141 488477
rect 101075 488412 101076 488476
rect 101140 488412 101141 488476
rect 101075 488411 101141 488412
rect 102363 488476 102429 488477
rect 102363 488412 102364 488476
rect 102428 488412 102429 488476
rect 102363 488411 102429 488412
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 475954 78914 488000
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 480454 83414 488000
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 484954 87914 488000
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 453454 92414 488000
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 457954 96914 488000
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 462454 101414 488000
rect 103286 487933 103346 489870
rect 104758 488477 104818 489870
rect 104755 488476 104821 488477
rect 104755 488412 104756 488476
rect 104820 488412 104821 488476
rect 104755 488411 104821 488412
rect 105310 488205 105370 489870
rect 105678 489870 105772 489930
rect 110462 489870 110532 489930
rect 115504 489930 115564 490106
rect 120536 489930 120596 490106
rect 125568 489930 125628 490106
rect 115504 489870 115674 489930
rect 120536 489870 120642 489930
rect 105678 488477 105738 489870
rect 105675 488476 105741 488477
rect 105675 488412 105676 488476
rect 105740 488412 105741 488476
rect 105675 488411 105741 488412
rect 110462 488205 110522 489870
rect 105307 488204 105373 488205
rect 105307 488140 105308 488204
rect 105372 488140 105373 488204
rect 105307 488139 105373 488140
rect 110459 488204 110525 488205
rect 110459 488140 110460 488204
rect 110524 488140 110525 488204
rect 110459 488139 110525 488140
rect 103283 487932 103349 487933
rect 103283 487868 103284 487932
rect 103348 487868 103349 487932
rect 103283 487867 103349 487868
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 466954 105914 488000
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 471454 110414 488000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 475954 114914 488000
rect 115614 487253 115674 489870
rect 115611 487252 115677 487253
rect 115611 487188 115612 487252
rect 115676 487188 115677 487252
rect 115611 487187 115677 487188
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 480454 119414 488000
rect 120582 487253 120642 489870
rect 125550 489870 125628 489930
rect 130464 489930 130524 490106
rect 135496 489930 135556 490106
rect 130464 489870 130578 489930
rect 120579 487252 120645 487253
rect 120579 487188 120580 487252
rect 120644 487188 120645 487252
rect 120579 487187 120645 487188
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 484954 123914 488000
rect 125550 487253 125610 489870
rect 125547 487252 125613 487253
rect 125547 487188 125548 487252
rect 125612 487188 125613 487252
rect 125547 487187 125613 487188
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 453454 128414 488000
rect 130518 487253 130578 489870
rect 135486 489870 135556 489930
rect 140528 489930 140588 490106
rect 140528 489870 140698 489930
rect 130515 487252 130581 487253
rect 130515 487188 130516 487252
rect 130580 487188 130581 487252
rect 130515 487187 130581 487188
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 457954 132914 488000
rect 135486 487253 135546 489870
rect 135483 487252 135549 487253
rect 135483 487188 135484 487252
rect 135548 487188 135549 487252
rect 135483 487187 135549 487188
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 462454 137414 488000
rect 140638 487253 140698 489870
rect 140635 487252 140701 487253
rect 140635 487188 140636 487252
rect 140700 487188 140701 487252
rect 140635 487187 140701 487188
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 466954 141914 488000
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 471454 146414 488000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 475954 150914 488000
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 480454 155414 488000
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 484954 159914 488000
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 453454 164414 488000
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 457954 168914 488000
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 462454 173414 488000
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 691292 191414 695898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 691292 195914 700398
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 691292 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 691292 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 691292 231914 700398
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 691292 258914 691398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 691292 263414 695898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 691292 267914 700398
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 190952 687454 191300 687486
rect 190952 687218 191008 687454
rect 191244 687218 191300 687454
rect 190952 687134 191300 687218
rect 190952 686898 191008 687134
rect 191244 686898 191300 687134
rect 190952 686866 191300 686898
rect 279760 687454 280108 687486
rect 279760 687218 279816 687454
rect 280052 687218 280108 687454
rect 279760 687134 280108 687218
rect 279760 686898 279816 687134
rect 280052 686898 280108 687134
rect 279760 686866 280108 686898
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 190272 655954 190620 655986
rect 190272 655718 190328 655954
rect 190564 655718 190620 655954
rect 190272 655634 190620 655718
rect 190272 655398 190328 655634
rect 190564 655398 190620 655634
rect 190272 655366 190620 655398
rect 280440 655954 280788 655986
rect 280440 655718 280496 655954
rect 280732 655718 280788 655954
rect 280440 655634 280788 655718
rect 280440 655398 280496 655634
rect 280732 655398 280788 655634
rect 280440 655366 280788 655398
rect 190952 651454 191300 651486
rect 190952 651218 191008 651454
rect 191244 651218 191300 651454
rect 190952 651134 191300 651218
rect 190952 650898 191008 651134
rect 191244 650898 191300 651134
rect 190952 650866 191300 650898
rect 279760 651454 280108 651486
rect 279760 651218 279816 651454
rect 280052 651218 280108 651454
rect 279760 651134 280108 651218
rect 279760 650898 279816 651134
rect 280052 650898 280108 651134
rect 279760 650866 280108 650898
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 190272 619954 190620 619986
rect 190272 619718 190328 619954
rect 190564 619718 190620 619954
rect 190272 619634 190620 619718
rect 190272 619398 190328 619634
rect 190564 619398 190620 619634
rect 190272 619366 190620 619398
rect 280440 619954 280788 619986
rect 280440 619718 280496 619954
rect 280732 619718 280788 619954
rect 280440 619634 280788 619718
rect 280440 619398 280496 619634
rect 280732 619398 280788 619634
rect 280440 619366 280788 619398
rect 190952 615454 191300 615486
rect 190952 615218 191008 615454
rect 191244 615218 191300 615454
rect 190952 615134 191300 615218
rect 190952 614898 191008 615134
rect 191244 614898 191300 615134
rect 190952 614866 191300 614898
rect 279760 615454 280108 615486
rect 279760 615218 279816 615454
rect 280052 615218 280108 615454
rect 279760 615134 280108 615218
rect 279760 614898 279816 615134
rect 280052 614898 280108 615134
rect 279760 614866 280108 614898
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 202928 599450 202988 600100
rect 202830 599390 202988 599450
rect 204288 599450 204348 600100
rect 205376 599450 205436 600100
rect 207688 599450 207748 600100
rect 208912 599450 208972 600100
rect 204288 599390 204362 599450
rect 205376 599390 205466 599450
rect 207688 599390 207858 599450
rect 202830 596461 202890 599390
rect 202827 596460 202893 596461
rect 202827 596396 202828 596460
rect 202892 596396 202893 596460
rect 202827 596395 202893 596396
rect 204302 596325 204362 599390
rect 205406 597141 205466 599390
rect 207798 597549 207858 599390
rect 208902 599390 208972 599450
rect 210000 599450 210060 600100
rect 211088 599450 211148 600100
rect 212312 599450 212372 600100
rect 213400 599450 213460 600100
rect 214760 599450 214820 600100
rect 215304 599450 215364 600100
rect 215712 599450 215772 600100
rect 220472 599450 220532 600100
rect 225504 599450 225564 600100
rect 210000 599390 210066 599450
rect 211088 599390 211170 599450
rect 212312 599390 212458 599450
rect 213400 599390 213562 599450
rect 214760 599390 214850 599450
rect 215304 599390 215402 599450
rect 208902 597549 208962 599390
rect 210006 597549 210066 599390
rect 211110 597549 211170 599390
rect 212398 597549 212458 599390
rect 213502 597549 213562 599390
rect 214790 597549 214850 599390
rect 215342 597549 215402 599390
rect 215710 599390 215772 599450
rect 219206 599390 220532 599450
rect 225462 599390 225564 599450
rect 230536 599450 230596 600100
rect 235568 599450 235628 600100
rect 240464 599450 240524 600100
rect 245496 599450 245556 600100
rect 250528 599450 250588 600100
rect 230536 599390 230674 599450
rect 235568 599390 235642 599450
rect 240464 599390 240610 599450
rect 245496 599390 245578 599450
rect 215710 597549 215770 599390
rect 207795 597548 207861 597549
rect 207795 597484 207796 597548
rect 207860 597484 207861 597548
rect 207795 597483 207861 597484
rect 208899 597548 208965 597549
rect 208899 597484 208900 597548
rect 208964 597484 208965 597548
rect 208899 597483 208965 597484
rect 210003 597548 210069 597549
rect 210003 597484 210004 597548
rect 210068 597484 210069 597548
rect 210003 597483 210069 597484
rect 211107 597548 211173 597549
rect 211107 597484 211108 597548
rect 211172 597484 211173 597548
rect 211107 597483 211173 597484
rect 212395 597548 212461 597549
rect 212395 597484 212396 597548
rect 212460 597484 212461 597548
rect 212395 597483 212461 597484
rect 213499 597548 213565 597549
rect 213499 597484 213500 597548
rect 213564 597484 213565 597548
rect 213499 597483 213565 597484
rect 214787 597548 214853 597549
rect 214787 597484 214788 597548
rect 214852 597484 214853 597548
rect 214787 597483 214853 597484
rect 215339 597548 215405 597549
rect 215339 597484 215340 597548
rect 215404 597484 215405 597548
rect 215339 597483 215405 597484
rect 215707 597548 215773 597549
rect 215707 597484 215708 597548
rect 215772 597484 215773 597548
rect 215707 597483 215773 597484
rect 205403 597140 205469 597141
rect 205403 597076 205404 597140
rect 205468 597076 205469 597140
rect 205403 597075 205469 597076
rect 219206 596325 219266 599390
rect 225462 597549 225522 599390
rect 225459 597548 225525 597549
rect 225459 597484 225460 597548
rect 225524 597484 225525 597548
rect 225459 597483 225525 597484
rect 230614 597277 230674 599390
rect 235582 597549 235642 599390
rect 235579 597548 235645 597549
rect 235579 597484 235580 597548
rect 235644 597484 235645 597548
rect 235579 597483 235645 597484
rect 230611 597276 230677 597277
rect 230611 597212 230612 597276
rect 230676 597212 230677 597276
rect 230611 597211 230677 597212
rect 240550 596869 240610 599390
rect 245518 597549 245578 599390
rect 250486 599390 250588 599450
rect 250486 597549 250546 599390
rect 245515 597548 245581 597549
rect 245515 597484 245516 597548
rect 245580 597484 245581 597548
rect 245515 597483 245581 597484
rect 250483 597548 250549 597549
rect 250483 597484 250484 597548
rect 250548 597484 250549 597548
rect 250483 597483 250549 597484
rect 240547 596868 240613 596869
rect 240547 596804 240548 596868
rect 240612 596804 240613 596868
rect 240547 596803 240613 596804
rect 204299 596324 204365 596325
rect 204299 596260 204300 596324
rect 204364 596260 204365 596324
rect 204299 596259 204365 596260
rect 219203 596324 219269 596325
rect 219203 596260 219204 596324
rect 219268 596260 219269 596324
rect 219203 596259 219269 596260
rect 282131 589932 282197 589933
rect 282131 589868 282132 589932
rect 282196 589868 282197 589932
rect 282131 589867 282197 589868
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 190272 547954 190620 547986
rect 190272 547718 190328 547954
rect 190564 547718 190620 547954
rect 190272 547634 190620 547718
rect 190272 547398 190328 547634
rect 190564 547398 190620 547634
rect 190272 547366 190620 547398
rect 280440 547954 280788 547986
rect 280440 547718 280496 547954
rect 280732 547718 280788 547954
rect 280440 547634 280788 547718
rect 280440 547398 280496 547634
rect 280732 547398 280788 547634
rect 280440 547366 280788 547398
rect 190952 543454 191300 543486
rect 190952 543218 191008 543454
rect 191244 543218 191300 543454
rect 190952 543134 191300 543218
rect 190952 542898 191008 543134
rect 191244 542898 191300 543134
rect 190952 542866 191300 542898
rect 279760 543454 280108 543486
rect 279760 543218 279816 543454
rect 280052 543218 280108 543454
rect 279760 543134 280108 543218
rect 279760 542898 279816 543134
rect 280052 542898 280108 543134
rect 279760 542866 280108 542898
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 190272 511954 190620 511986
rect 190272 511718 190328 511954
rect 190564 511718 190620 511954
rect 190272 511634 190620 511718
rect 190272 511398 190328 511634
rect 190564 511398 190620 511634
rect 190272 511366 190620 511398
rect 280440 511954 280788 511986
rect 280440 511718 280496 511954
rect 280732 511718 280788 511954
rect 280440 511634 280788 511718
rect 280440 511398 280496 511634
rect 280732 511398 280788 511634
rect 280440 511366 280788 511398
rect 190952 507454 191300 507486
rect 190952 507218 191008 507454
rect 191244 507218 191300 507454
rect 190952 507134 191300 507218
rect 190952 506898 191008 507134
rect 191244 506898 191300 507134
rect 190952 506866 191300 506898
rect 279760 507454 280108 507486
rect 279760 507218 279816 507454
rect 280052 507218 280108 507454
rect 279760 507134 280108 507218
rect 279760 506898 279816 507134
rect 280052 506898 280108 507134
rect 279760 506866 280108 506898
rect 202928 489930 202988 490106
rect 204288 489930 204348 490106
rect 205376 489930 205436 490106
rect 207688 489930 207748 490106
rect 208912 489930 208972 490106
rect 202928 489870 203074 489930
rect 204288 489870 204362 489930
rect 205376 489870 205466 489930
rect 203014 488205 203074 489870
rect 204302 488477 204362 489870
rect 204299 488476 204365 488477
rect 204299 488412 204300 488476
rect 204364 488412 204365 488476
rect 204299 488411 204365 488412
rect 203011 488204 203077 488205
rect 203011 488140 203012 488204
rect 203076 488140 203077 488204
rect 203011 488139 203077 488140
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 480454 191414 488000
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 484954 195914 488000
rect 203014 487253 203074 488139
rect 205406 487253 205466 489870
rect 207614 489870 207748 489930
rect 208902 489870 208972 489930
rect 210000 489930 210060 490106
rect 211088 489930 211148 490106
rect 212312 489930 212372 490106
rect 210000 489870 210066 489930
rect 211088 489870 211170 489930
rect 207614 487253 207674 489870
rect 208902 487933 208962 489870
rect 208899 487932 208965 487933
rect 208899 487868 208900 487932
rect 208964 487868 208965 487932
rect 208899 487867 208965 487868
rect 210006 487253 210066 489870
rect 211110 488341 211170 489870
rect 212214 489870 212372 489930
rect 213400 489930 213460 490106
rect 214760 489930 214820 490106
rect 215304 489930 215364 490106
rect 215712 489930 215772 490106
rect 213400 489870 213562 489930
rect 214760 489870 214850 489930
rect 215304 489870 215402 489930
rect 211107 488340 211173 488341
rect 211107 488276 211108 488340
rect 211172 488276 211173 488340
rect 211107 488275 211173 488276
rect 212214 487525 212274 489870
rect 213502 488341 213562 489870
rect 214790 488477 214850 489870
rect 214787 488476 214853 488477
rect 214787 488412 214788 488476
rect 214852 488412 214853 488476
rect 214787 488411 214853 488412
rect 213499 488340 213565 488341
rect 213499 488276 213500 488340
rect 213564 488276 213565 488340
rect 213499 488275 213565 488276
rect 212211 487524 212277 487525
rect 212211 487460 212212 487524
rect 212276 487460 212277 487524
rect 212211 487459 212277 487460
rect 215342 487253 215402 489870
rect 215710 489870 215772 489930
rect 220472 489930 220532 490106
rect 225504 489930 225564 490106
rect 220472 489870 220554 489930
rect 215710 488341 215770 489870
rect 215707 488340 215773 488341
rect 215707 488276 215708 488340
rect 215772 488276 215773 488340
rect 215707 488275 215773 488276
rect 220494 487253 220554 489870
rect 225462 489870 225564 489930
rect 230536 489930 230596 490106
rect 235568 489930 235628 490106
rect 240464 489930 240524 490106
rect 245496 489930 245556 490106
rect 250528 489930 250588 490106
rect 230536 489870 230674 489930
rect 235568 489870 235642 489930
rect 240464 489870 240610 489930
rect 245496 489870 245578 489930
rect 225462 487253 225522 489870
rect 230614 487253 230674 489870
rect 203011 487252 203077 487253
rect 203011 487188 203012 487252
rect 203076 487188 203077 487252
rect 203011 487187 203077 487188
rect 205403 487252 205469 487253
rect 205403 487188 205404 487252
rect 205468 487188 205469 487252
rect 205403 487187 205469 487188
rect 207611 487252 207677 487253
rect 207611 487188 207612 487252
rect 207676 487188 207677 487252
rect 207611 487187 207677 487188
rect 210003 487252 210069 487253
rect 210003 487188 210004 487252
rect 210068 487188 210069 487252
rect 210003 487187 210069 487188
rect 215339 487252 215405 487253
rect 215339 487188 215340 487252
rect 215404 487188 215405 487252
rect 215339 487187 215405 487188
rect 220491 487252 220557 487253
rect 220491 487188 220492 487252
rect 220556 487188 220557 487252
rect 220491 487187 220557 487188
rect 225459 487252 225525 487253
rect 225459 487188 225460 487252
rect 225524 487188 225525 487252
rect 225459 487187 225525 487188
rect 230611 487252 230677 487253
rect 230611 487188 230612 487252
rect 230676 487188 230677 487252
rect 230611 487187 230677 487188
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 231294 484954 231914 488000
rect 235582 487253 235642 489870
rect 240550 487253 240610 489870
rect 245518 487253 245578 489870
rect 250486 489870 250588 489930
rect 250486 487253 250546 489870
rect 235579 487252 235645 487253
rect 235579 487188 235580 487252
rect 235644 487188 235645 487252
rect 235579 487187 235645 487188
rect 240547 487252 240613 487253
rect 240547 487188 240548 487252
rect 240612 487188 240613 487252
rect 240547 487187 240613 487188
rect 245515 487252 245581 487253
rect 245515 487188 245516 487252
rect 245580 487188 245581 487252
rect 245515 487187 245581 487188
rect 250483 487252 250549 487253
rect 250483 487188 250484 487252
rect 250548 487188 250549 487252
rect 250483 487187 250549 487188
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 446000 231914 448398
rect 267294 484954 267914 488000
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 258579 446588 258645 446589
rect 258579 446524 258580 446588
rect 258644 446524 258645 446588
rect 258579 446523 258645 446524
rect 209635 444140 209701 444141
rect 209635 444076 209636 444140
rect 209700 444076 209701 444140
rect 209635 444075 209701 444076
rect 210739 444140 210805 444141
rect 210739 444076 210740 444140
rect 210804 444076 210805 444140
rect 210739 444075 210805 444076
rect 238155 444140 238221 444141
rect 238155 444076 238156 444140
rect 238220 444076 238221 444140
rect 238155 444075 238221 444076
rect 256371 444140 256437 444141
rect 256371 444076 256372 444140
rect 256436 444076 256437 444140
rect 256371 444075 256437 444076
rect 203379 443052 203445 443053
rect 203379 442988 203380 443052
rect 203444 442988 203445 443052
rect 203379 442987 203445 442988
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 381454 200414 398000
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 203382 292637 203442 442987
rect 209638 442237 209698 444075
rect 210742 442373 210802 444075
rect 220123 443732 220189 443733
rect 220123 443668 220124 443732
rect 220188 443668 220189 443732
rect 220123 443667 220189 443668
rect 220126 443053 220186 443667
rect 220123 443052 220189 443053
rect 220123 442988 220124 443052
rect 220188 442988 220189 443052
rect 220123 442987 220189 442988
rect 238158 442509 238218 444075
rect 245515 444004 245581 444005
rect 245515 443940 245516 444004
rect 245580 443940 245581 444004
rect 245515 443939 245581 443940
rect 251035 444004 251101 444005
rect 251035 443940 251036 444004
rect 251100 443940 251101 444004
rect 251035 443939 251101 443940
rect 245518 442645 245578 443939
rect 251038 442781 251098 443939
rect 251035 442780 251101 442781
rect 251035 442716 251036 442780
rect 251100 442716 251101 442780
rect 251035 442715 251101 442716
rect 245515 442644 245581 442645
rect 245515 442580 245516 442644
rect 245580 442580 245581 442644
rect 245515 442579 245581 442580
rect 238155 442508 238221 442509
rect 238155 442444 238156 442508
rect 238220 442444 238221 442508
rect 238155 442443 238221 442444
rect 210739 442372 210805 442373
rect 210739 442308 210740 442372
rect 210804 442308 210805 442372
rect 210739 442307 210805 442308
rect 209635 442236 209701 442237
rect 209635 442172 209636 442236
rect 209700 442172 209701 442236
rect 209635 442171 209701 442172
rect 256374 441693 256434 444075
rect 256371 441692 256437 441693
rect 256371 441628 256372 441692
rect 256436 441628 256437 441692
rect 256371 441627 256437 441628
rect 219568 439954 219888 439986
rect 219568 439718 219610 439954
rect 219846 439718 219888 439954
rect 219568 439634 219888 439718
rect 219568 439398 219610 439634
rect 219846 439398 219888 439634
rect 219568 439366 219888 439398
rect 250288 439954 250608 439986
rect 250288 439718 250330 439954
rect 250566 439718 250608 439954
rect 250288 439634 250608 439718
rect 250288 439398 250330 439634
rect 250566 439398 250608 439634
rect 250288 439366 250608 439398
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 219568 403954 219888 403986
rect 219568 403718 219610 403954
rect 219846 403718 219888 403954
rect 219568 403634 219888 403718
rect 219568 403398 219610 403634
rect 219846 403398 219888 403634
rect 219568 403366 219888 403398
rect 250288 403954 250608 403986
rect 250288 403718 250330 403954
rect 250566 403718 250608 403954
rect 250288 403634 250608 403718
rect 250288 403398 250330 403634
rect 250566 403398 250608 403634
rect 250288 403366 250608 403398
rect 252875 399940 252941 399941
rect 252875 399876 252876 399940
rect 252940 399876 252941 399940
rect 252875 399875 252941 399876
rect 252691 399260 252757 399261
rect 252691 399196 252692 399260
rect 252756 399196 252757 399260
rect 252691 399195 252757 399196
rect 252694 398853 252754 399195
rect 250299 398852 250365 398853
rect 250299 398788 250300 398852
rect 250364 398788 250365 398852
rect 250299 398787 250365 398788
rect 252691 398852 252757 398853
rect 252691 398788 252692 398852
rect 252756 398788 252757 398852
rect 252691 398787 252757 398788
rect 214603 398716 214669 398717
rect 214603 398652 214604 398716
rect 214668 398652 214669 398716
rect 214603 398651 214669 398652
rect 205587 398444 205653 398445
rect 205587 398380 205588 398444
rect 205652 398380 205653 398444
rect 205587 398379 205653 398380
rect 205590 398173 205650 398379
rect 211291 398308 211357 398309
rect 211291 398244 211292 398308
rect 211356 398244 211357 398308
rect 211291 398243 211357 398244
rect 205587 398172 205653 398173
rect 205587 398108 205588 398172
rect 205652 398108 205653 398172
rect 205587 398107 205653 398108
rect 204294 385954 204914 398000
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 203379 292636 203445 292637
rect 203379 292572 203380 292636
rect 203444 292572 203445 292636
rect 203379 292571 203445 292572
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 390454 209414 398000
rect 211294 397762 211354 398243
rect 211110 397702 211354 397762
rect 211659 397764 211725 397765
rect 209819 397628 209885 397629
rect 209819 397564 209820 397628
rect 209884 397564 209885 397628
rect 209819 397563 209885 397564
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 209822 8941 209882 397563
rect 210003 397492 210069 397493
rect 210003 397428 210004 397492
rect 210068 397428 210069 397492
rect 210003 397427 210069 397428
rect 210006 9077 210066 397427
rect 211110 392597 211170 397702
rect 211659 397700 211660 397764
rect 211724 397700 211725 397764
rect 211659 397699 211725 397700
rect 212763 397764 212829 397765
rect 212763 397700 212764 397764
rect 212828 397700 212829 397764
rect 212763 397699 212829 397700
rect 211291 397628 211357 397629
rect 211291 397564 211292 397628
rect 211356 397564 211357 397628
rect 211291 397563 211357 397564
rect 211107 392596 211173 392597
rect 211107 392532 211108 392596
rect 211172 392532 211173 392596
rect 211107 392531 211173 392532
rect 211294 11661 211354 397563
rect 211475 397492 211541 397493
rect 211475 397428 211476 397492
rect 211540 397428 211541 397492
rect 211475 397427 211541 397428
rect 211478 13157 211538 397427
rect 211475 13156 211541 13157
rect 211475 13092 211476 13156
rect 211540 13092 211541 13156
rect 211475 13091 211541 13092
rect 211291 11660 211357 11661
rect 211291 11596 211292 11660
rect 211356 11596 211357 11660
rect 211291 11595 211357 11596
rect 211662 9213 211722 397699
rect 212579 397492 212645 397493
rect 212579 397428 212580 397492
rect 212644 397428 212645 397492
rect 212579 397427 212645 397428
rect 212582 11797 212642 397427
rect 212766 395317 212826 397699
rect 212763 395316 212829 395317
rect 212763 395252 212764 395316
rect 212828 395252 212829 395316
rect 212763 395251 212829 395252
rect 213294 394954 213914 398000
rect 214051 397764 214117 397765
rect 214051 397700 214052 397764
rect 214116 397700 214117 397764
rect 214051 397699 214117 397700
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 212579 11796 212645 11797
rect 212579 11732 212580 11796
rect 212644 11732 212645 11796
rect 212579 11731 212645 11732
rect 211659 9212 211725 9213
rect 211659 9148 211660 9212
rect 211724 9148 211725 9212
rect 211659 9147 211725 9148
rect 210003 9076 210069 9077
rect 210003 9012 210004 9076
rect 210068 9012 210069 9076
rect 210003 9011 210069 9012
rect 209819 8940 209885 8941
rect 209819 8876 209820 8940
rect 209884 8876 209885 8940
rect 209819 8875 209885 8876
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 -7066 213914 34398
rect 214054 7581 214114 397699
rect 214419 397628 214485 397629
rect 214419 397564 214420 397628
rect 214484 397564 214485 397628
rect 214419 397563 214485 397564
rect 214235 397492 214301 397493
rect 214235 397428 214236 397492
rect 214300 397428 214301 397492
rect 214235 397427 214301 397428
rect 214238 11933 214298 397427
rect 214422 14517 214482 397563
rect 214606 395453 214666 398651
rect 228587 398580 228653 398581
rect 228587 398516 228588 398580
rect 228652 398516 228653 398580
rect 228587 398515 228653 398516
rect 216627 397900 216693 397901
rect 216627 397836 216628 397900
rect 216692 397836 216693 397900
rect 216627 397835 216693 397836
rect 215339 397764 215405 397765
rect 215339 397700 215340 397764
rect 215404 397700 215405 397764
rect 215339 397699 215405 397700
rect 215342 395589 215402 397699
rect 215707 397628 215773 397629
rect 215707 397564 215708 397628
rect 215772 397564 215773 397628
rect 215707 397563 215773 397564
rect 215523 397492 215589 397493
rect 215523 397428 215524 397492
rect 215588 397428 215589 397492
rect 215523 397427 215589 397428
rect 215339 395588 215405 395589
rect 215339 395524 215340 395588
rect 215404 395524 215405 395588
rect 215339 395523 215405 395524
rect 214603 395452 214669 395453
rect 214603 395388 214604 395452
rect 214668 395388 214669 395452
rect 214603 395387 214669 395388
rect 215526 177309 215586 397427
rect 215523 177308 215589 177309
rect 215523 177244 215524 177308
rect 215588 177244 215589 177308
rect 215523 177243 215589 177244
rect 214419 14516 214485 14517
rect 214419 14452 214420 14516
rect 214484 14452 214485 14516
rect 214419 14451 214485 14452
rect 215710 13021 215770 397563
rect 215707 13020 215773 13021
rect 215707 12956 215708 13020
rect 215772 12956 215773 13020
rect 215707 12955 215773 12956
rect 214235 11932 214301 11933
rect 214235 11868 214236 11932
rect 214300 11868 214301 11932
rect 214235 11867 214301 11868
rect 216630 10437 216690 397835
rect 216995 397764 217061 397765
rect 216995 397700 216996 397764
rect 217060 397700 217061 397764
rect 216995 397699 217061 397700
rect 216811 397492 216877 397493
rect 216811 397428 216812 397492
rect 216876 397428 216877 397492
rect 216811 397427 216877 397428
rect 216627 10436 216693 10437
rect 216627 10372 216628 10436
rect 216692 10372 216693 10436
rect 216627 10371 216693 10372
rect 216814 10301 216874 397427
rect 216998 14653 217058 397699
rect 217179 397628 217245 397629
rect 217179 397564 217180 397628
rect 217244 397564 217245 397628
rect 217179 397563 217245 397564
rect 217182 353973 217242 397563
rect 217794 363454 218414 398000
rect 218835 397628 218901 397629
rect 218835 397564 218836 397628
rect 218900 397564 218901 397628
rect 218835 397563 218901 397564
rect 219571 397628 219637 397629
rect 219571 397564 219572 397628
rect 219636 397564 219637 397628
rect 219571 397563 219637 397564
rect 220859 397628 220925 397629
rect 220859 397564 220860 397628
rect 220924 397564 220925 397628
rect 220859 397563 220925 397564
rect 221411 397628 221477 397629
rect 221411 397564 221412 397628
rect 221476 397564 221477 397628
rect 221411 397563 221477 397564
rect 218651 397492 218717 397493
rect 218651 397428 218652 397492
rect 218716 397428 218717 397492
rect 218651 397427 218717 397428
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217179 353972 217245 353973
rect 217179 353908 217180 353972
rect 217244 353908 217245 353972
rect 217179 353907 217245 353908
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 216995 14652 217061 14653
rect 216995 14588 216996 14652
rect 217060 14588 217061 14652
rect 216995 14587 217061 14588
rect 216811 10300 216877 10301
rect 216811 10236 216812 10300
rect 216876 10236 216877 10300
rect 216811 10235 216877 10236
rect 214051 7580 214117 7581
rect 214051 7516 214052 7580
rect 214116 7516 214117 7580
rect 214051 7515 214117 7516
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 3454 218414 38898
rect 218654 15877 218714 397427
rect 218838 354109 218898 397563
rect 219387 397492 219453 397493
rect 219387 397428 219388 397492
rect 219452 397428 219453 397492
rect 219387 397427 219453 397428
rect 219390 389190 219450 397427
rect 219206 389130 219450 389190
rect 218835 354108 218901 354109
rect 218835 354044 218836 354108
rect 218900 354044 218901 354108
rect 218835 354043 218901 354044
rect 218651 15876 218717 15877
rect 218651 15812 218652 15876
rect 218716 15812 218717 15876
rect 218651 15811 218717 15812
rect 219206 10573 219266 389130
rect 219574 12069 219634 397563
rect 219755 397492 219821 397493
rect 219755 397428 219756 397492
rect 219820 397428 219821 397492
rect 219755 397427 219821 397428
rect 219758 177445 219818 397427
rect 220862 393957 220922 397563
rect 221043 397492 221109 397493
rect 221043 397428 221044 397492
rect 221108 397428 221109 397492
rect 221043 397427 221109 397428
rect 221227 397492 221293 397493
rect 221227 397428 221228 397492
rect 221292 397428 221293 397492
rect 221227 397427 221293 397428
rect 220859 393956 220925 393957
rect 220859 393892 220860 393956
rect 220924 393892 220925 393956
rect 220859 393891 220925 393892
rect 219755 177444 219821 177445
rect 219755 177380 219756 177444
rect 219820 177380 219821 177444
rect 219755 177379 219821 177380
rect 219571 12068 219637 12069
rect 219571 12004 219572 12068
rect 219636 12004 219637 12068
rect 219571 12003 219637 12004
rect 219203 10572 219269 10573
rect 219203 10508 219204 10572
rect 219268 10508 219269 10572
rect 219203 10507 219269 10508
rect 221046 7717 221106 397427
rect 221230 394093 221290 397427
rect 221227 394092 221293 394093
rect 221227 394028 221228 394092
rect 221292 394028 221293 394092
rect 221227 394027 221293 394028
rect 221414 7853 221474 397563
rect 222147 397492 222213 397493
rect 222147 397428 222148 397492
rect 222212 397428 222213 397492
rect 222147 397427 222213 397428
rect 222150 394229 222210 397427
rect 222147 394228 222213 394229
rect 222147 394164 222148 394228
rect 222212 394164 222213 394228
rect 222147 394163 222213 394164
rect 222294 367954 222914 398000
rect 223987 397900 224053 397901
rect 223987 397836 223988 397900
rect 224052 397836 224053 397900
rect 223987 397835 224053 397836
rect 224907 397900 224973 397901
rect 224907 397836 224908 397900
rect 224972 397836 224973 397900
rect 224907 397835 224973 397836
rect 223067 397764 223133 397765
rect 223067 397700 223068 397764
rect 223132 397700 223133 397764
rect 223067 397699 223133 397700
rect 223070 392733 223130 397699
rect 223619 397628 223685 397629
rect 223619 397564 223620 397628
rect 223684 397564 223685 397628
rect 223619 397563 223685 397564
rect 223067 392732 223133 392733
rect 223067 392668 223068 392732
rect 223132 392668 223133 392732
rect 223067 392667 223133 392668
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 221411 7852 221477 7853
rect 221411 7788 221412 7852
rect 221476 7788 221477 7852
rect 221411 7787 221477 7788
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 221043 7716 221109 7717
rect 221043 7652 221044 7716
rect 221108 7652 221109 7716
rect 221043 7651 221109 7652
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 223622 3365 223682 397563
rect 223803 397492 223869 397493
rect 223803 397428 223804 397492
rect 223868 397428 223869 397492
rect 223803 397427 223869 397428
rect 223806 6221 223866 397427
rect 223990 16013 224050 397835
rect 224171 397764 224237 397765
rect 224171 397700 224172 397764
rect 224236 397700 224237 397764
rect 224910 397762 224970 397835
rect 224171 397699 224237 397700
rect 224726 397702 224970 397762
rect 225275 397764 225341 397765
rect 224174 177581 224234 397699
rect 224726 389190 224786 397702
rect 225275 397700 225276 397764
rect 225340 397700 225341 397764
rect 225275 397699 225341 397700
rect 225091 397492 225157 397493
rect 225091 397428 225092 397492
rect 225156 397428 225157 397492
rect 225091 397427 225157 397428
rect 224726 389130 224970 389190
rect 224171 177580 224237 177581
rect 224171 177516 224172 177580
rect 224236 177516 224237 177580
rect 224171 177515 224237 177516
rect 223987 16012 224053 16013
rect 223987 15948 223988 16012
rect 224052 15948 224053 16012
rect 223987 15947 224053 15948
rect 224910 6357 224970 389130
rect 225094 46205 225154 397427
rect 225278 178669 225338 397699
rect 225459 397628 225525 397629
rect 225459 397564 225460 397628
rect 225524 397564 225525 397628
rect 225459 397563 225525 397564
rect 226563 397628 226629 397629
rect 226563 397564 226564 397628
rect 226628 397564 226629 397628
rect 226563 397563 226629 397564
rect 225462 352613 225522 397563
rect 225459 352612 225525 352613
rect 225459 352548 225460 352612
rect 225524 352548 225525 352612
rect 225459 352547 225525 352548
rect 225275 178668 225341 178669
rect 225275 178604 225276 178668
rect 225340 178604 225341 178668
rect 225275 178603 225341 178604
rect 225091 46204 225157 46205
rect 225091 46140 225092 46204
rect 225156 46140 225157 46204
rect 225091 46139 225157 46140
rect 224907 6356 224973 6357
rect 224907 6292 224908 6356
rect 224972 6292 224973 6356
rect 224907 6291 224973 6292
rect 223803 6220 223869 6221
rect 223803 6156 223804 6220
rect 223868 6156 223869 6220
rect 223803 6155 223869 6156
rect 226566 3909 226626 397563
rect 226794 372454 227414 398000
rect 228403 397764 228469 397765
rect 228403 397700 228404 397764
rect 228468 397700 228469 397764
rect 228403 397699 228469 397700
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226563 3908 226629 3909
rect 226563 3844 226564 3908
rect 226628 3844 226629 3908
rect 226563 3843 226629 3844
rect 223619 3364 223685 3365
rect 223619 3300 223620 3364
rect 223684 3300 223685 3364
rect 223619 3299 223685 3300
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 -2266 227414 11898
rect 228406 6357 228466 397699
rect 228403 6356 228469 6357
rect 228403 6292 228404 6356
rect 228468 6292 228469 6356
rect 228403 6291 228469 6292
rect 228590 4045 228650 398515
rect 246987 398308 247053 398309
rect 246987 398244 246988 398308
rect 247052 398244 247053 398308
rect 246987 398243 247053 398244
rect 230427 398036 230493 398037
rect 230427 397972 230428 398036
rect 230492 397972 230493 398036
rect 233187 398036 233253 398037
rect 230427 397971 230493 397972
rect 228771 397900 228837 397901
rect 228771 397836 228772 397900
rect 228836 397836 228837 397900
rect 228771 397835 228837 397836
rect 228587 4044 228653 4045
rect 228587 3980 228588 4044
rect 228652 3980 228653 4044
rect 228587 3979 228653 3980
rect 228774 3501 228834 397835
rect 230059 397764 230125 397765
rect 230059 397700 230060 397764
rect 230124 397700 230125 397764
rect 230059 397699 230125 397700
rect 229875 397628 229941 397629
rect 229875 397564 229876 397628
rect 229940 397564 229941 397628
rect 229875 397563 229941 397564
rect 228955 397492 229021 397493
rect 228955 397428 228956 397492
rect 229020 397428 229021 397492
rect 228955 397427 229021 397428
rect 228958 3637 229018 397427
rect 229878 5133 229938 397563
rect 230062 5541 230122 397699
rect 230243 397492 230309 397493
rect 230243 397428 230244 397492
rect 230308 397428 230309 397492
rect 230243 397427 230309 397428
rect 230059 5540 230125 5541
rect 230059 5476 230060 5540
rect 230124 5476 230125 5540
rect 230059 5475 230125 5476
rect 229875 5132 229941 5133
rect 229875 5068 229876 5132
rect 229940 5068 229941 5132
rect 229875 5067 229941 5068
rect 228955 3636 229021 3637
rect 228955 3572 228956 3636
rect 229020 3572 229021 3636
rect 228955 3571 229021 3572
rect 228771 3500 228837 3501
rect 228771 3436 228772 3500
rect 228836 3436 228837 3500
rect 228771 3435 228837 3436
rect 230246 3365 230306 397427
rect 230430 395725 230490 397971
rect 230611 397764 230677 397765
rect 230611 397700 230612 397764
rect 230676 397700 230677 397764
rect 230611 397699 230677 397700
rect 230427 395724 230493 395725
rect 230427 395660 230428 395724
rect 230492 395660 230493 395724
rect 230427 395659 230493 395660
rect 230614 354381 230674 397699
rect 230795 397628 230861 397629
rect 230795 397564 230796 397628
rect 230860 397564 230861 397628
rect 230795 397563 230861 397564
rect 230611 354380 230677 354381
rect 230611 354316 230612 354380
rect 230676 354316 230677 354380
rect 230611 354315 230677 354316
rect 230798 6765 230858 397563
rect 230979 397492 231045 397493
rect 230979 397428 230980 397492
rect 231044 397428 231045 397492
rect 230979 397427 231045 397428
rect 230795 6764 230861 6765
rect 230795 6700 230796 6764
rect 230860 6700 230861 6764
rect 230795 6699 230861 6700
rect 230243 3364 230309 3365
rect 230243 3300 230244 3364
rect 230308 3300 230309 3364
rect 230243 3299 230309 3300
rect 230982 3229 231042 397427
rect 231294 376954 231914 398000
rect 233187 397972 233188 398036
rect 233252 397972 233253 398036
rect 233187 397971 233253 397972
rect 232819 397764 232885 397765
rect 232819 397700 232820 397764
rect 232884 397700 232885 397764
rect 232819 397699 232885 397700
rect 232635 397628 232701 397629
rect 232635 397564 232636 397628
rect 232700 397564 232701 397628
rect 232635 397563 232701 397564
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 232638 18869 232698 397563
rect 232635 18868 232701 18869
rect 232635 18804 232636 18868
rect 232700 18804 232701 18868
rect 232635 18803 232701 18804
rect 232822 18733 232882 397699
rect 233003 397492 233069 397493
rect 233003 397428 233004 397492
rect 233068 397428 233069 397492
rect 233003 397427 233069 397428
rect 232819 18732 232885 18733
rect 232819 18668 232820 18732
rect 232884 18668 232885 18732
rect 232819 18667 232885 18668
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 230979 3228 231045 3229
rect 230979 3164 230980 3228
rect 231044 3164 231045 3228
rect 230979 3163 231045 3164
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 -3226 231914 16398
rect 233006 6629 233066 397427
rect 233190 395589 233250 397971
rect 233923 397764 233989 397765
rect 233923 397700 233924 397764
rect 233988 397700 233989 397764
rect 233923 397699 233989 397700
rect 235211 397764 235277 397765
rect 235211 397700 235212 397764
rect 235276 397700 235277 397764
rect 235211 397699 235277 397700
rect 233187 395588 233253 395589
rect 233187 395524 233188 395588
rect 233252 395524 233253 395588
rect 233187 395523 233253 395524
rect 233926 7717 233986 397699
rect 234107 397628 234173 397629
rect 234107 397564 234108 397628
rect 234172 397564 234173 397628
rect 234107 397563 234173 397564
rect 234110 25533 234170 397563
rect 234291 397492 234357 397493
rect 234291 397428 234292 397492
rect 234356 397428 234357 397492
rect 234291 397427 234357 397428
rect 234107 25532 234173 25533
rect 234107 25468 234108 25532
rect 234172 25468 234173 25532
rect 234107 25467 234173 25468
rect 234294 18597 234354 397427
rect 235214 83469 235274 397699
rect 235395 397628 235461 397629
rect 235395 397564 235396 397628
rect 235460 397564 235461 397628
rect 235395 397563 235461 397564
rect 235211 83468 235277 83469
rect 235211 83404 235212 83468
rect 235276 83404 235277 83468
rect 235211 83403 235277 83404
rect 234291 18596 234357 18597
rect 234291 18532 234292 18596
rect 234356 18532 234357 18596
rect 234291 18531 234357 18532
rect 235398 9077 235458 397563
rect 235579 397492 235645 397493
rect 235579 397428 235580 397492
rect 235644 397428 235645 397492
rect 235579 397427 235645 397428
rect 235395 9076 235461 9077
rect 235395 9012 235396 9076
rect 235460 9012 235461 9076
rect 235395 9011 235461 9012
rect 233923 7716 233989 7717
rect 233923 7652 233924 7716
rect 233988 7652 233989 7716
rect 233923 7651 233989 7652
rect 235582 7581 235642 397427
rect 235794 381454 236414 398000
rect 236867 397764 236933 397765
rect 236867 397700 236868 397764
rect 236932 397700 236933 397764
rect 236867 397699 236933 397700
rect 238155 397764 238221 397765
rect 238155 397700 238156 397764
rect 238220 397700 238221 397764
rect 238155 397699 238221 397700
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 236870 27029 236930 397699
rect 237051 397628 237117 397629
rect 237051 397564 237052 397628
rect 237116 397564 237117 397628
rect 237051 397563 237117 397564
rect 236867 27028 236933 27029
rect 236867 26964 236868 27028
rect 236932 26964 236933 27028
rect 236867 26963 236933 26964
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235579 7580 235645 7581
rect 235579 7516 235580 7580
rect 235644 7516 235645 7580
rect 235579 7515 235645 7516
rect 233003 6628 233069 6629
rect 233003 6564 233004 6628
rect 233068 6564 233069 6628
rect 233003 6563 233069 6564
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 -4186 236414 20898
rect 237054 19957 237114 397563
rect 237235 397492 237301 397493
rect 237235 397428 237236 397492
rect 237300 397428 237301 397492
rect 237235 397427 237301 397428
rect 237051 19956 237117 19957
rect 237051 19892 237052 19956
rect 237116 19892 237117 19956
rect 237051 19891 237117 19892
rect 237238 6493 237298 397427
rect 238158 352885 238218 397699
rect 238339 397628 238405 397629
rect 238339 397564 238340 397628
rect 238404 397564 238405 397628
rect 238339 397563 238405 397564
rect 239811 397628 239877 397629
rect 239811 397564 239812 397628
rect 239876 397564 239877 397628
rect 239811 397563 239877 397564
rect 238155 352884 238221 352885
rect 238155 352820 238156 352884
rect 238220 352820 238221 352884
rect 238155 352819 238221 352820
rect 238342 26893 238402 397563
rect 238523 397492 238589 397493
rect 238523 397428 238524 397492
rect 238588 397428 238589 397492
rect 238523 397427 238589 397428
rect 239627 397492 239693 397493
rect 239627 397428 239628 397492
rect 239692 397428 239693 397492
rect 239627 397427 239693 397428
rect 238339 26892 238405 26893
rect 238339 26828 238340 26892
rect 238404 26828 238405 26892
rect 238339 26827 238405 26828
rect 238526 8941 238586 397427
rect 239630 21725 239690 397427
rect 239627 21724 239693 21725
rect 239627 21660 239628 21724
rect 239692 21660 239693 21724
rect 239627 21659 239693 21660
rect 239814 21589 239874 397563
rect 239995 397492 240061 397493
rect 239995 397428 239996 397492
rect 240060 397428 240061 397492
rect 239995 397427 240061 397428
rect 239811 21588 239877 21589
rect 239811 21524 239812 21588
rect 239876 21524 239877 21588
rect 239811 21523 239877 21524
rect 239998 10573 240058 397427
rect 240294 385954 240914 398000
rect 242387 397900 242453 397901
rect 242387 397836 242388 397900
rect 242452 397836 242453 397900
rect 242387 397835 242453 397836
rect 242203 397764 242269 397765
rect 242203 397700 242204 397764
rect 242268 397700 242269 397764
rect 242203 397699 242269 397700
rect 241283 397492 241349 397493
rect 241283 397428 241284 397492
rect 241348 397428 241349 397492
rect 241283 397427 241349 397428
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 241286 351117 241346 397427
rect 241283 351116 241349 351117
rect 241283 351052 241284 351116
rect 241348 351052 241349 351116
rect 241283 351051 241349 351052
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 239995 10572 240061 10573
rect 239995 10508 239996 10572
rect 240060 10508 240061 10572
rect 239995 10507 240061 10508
rect 238523 8940 238589 8941
rect 238523 8876 238524 8940
rect 238588 8876 238589 8940
rect 238523 8875 238589 8876
rect 237235 6492 237301 6493
rect 237235 6428 237236 6492
rect 237300 6428 237301 6492
rect 237235 6427 237301 6428
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 -5146 240914 25398
rect 242206 21453 242266 397699
rect 242203 21452 242269 21453
rect 242203 21388 242204 21452
rect 242268 21388 242269 21452
rect 242203 21387 242269 21388
rect 242390 21317 242450 397835
rect 243675 397764 243741 397765
rect 243675 397700 243676 397764
rect 243740 397700 243741 397764
rect 243675 397699 243741 397700
rect 242755 397628 242821 397629
rect 242755 397564 242756 397628
rect 242820 397564 242821 397628
rect 242755 397563 242821 397564
rect 242571 397492 242637 397493
rect 242571 397428 242572 397492
rect 242636 397428 242637 397492
rect 242571 397427 242637 397428
rect 242387 21316 242453 21317
rect 242387 21252 242388 21316
rect 242452 21252 242453 21316
rect 242387 21251 242453 21252
rect 242574 10301 242634 397427
rect 242758 10437 242818 397563
rect 243678 177309 243738 397699
rect 244043 397628 244109 397629
rect 244043 397564 244044 397628
rect 244108 397564 244109 397628
rect 244043 397563 244109 397564
rect 243859 397492 243925 397493
rect 243859 397428 243860 397492
rect 243924 397428 243925 397492
rect 243859 397427 243925 397428
rect 243675 177308 243741 177309
rect 243675 177244 243676 177308
rect 243740 177244 243741 177308
rect 243675 177243 243741 177244
rect 243862 16285 243922 397427
rect 243859 16284 243925 16285
rect 243859 16220 243860 16284
rect 243924 16220 243925 16284
rect 243859 16219 243925 16220
rect 244046 11797 244106 397563
rect 244794 390454 245414 398000
rect 246435 397764 246501 397765
rect 246435 397700 246436 397764
rect 246500 397700 246501 397764
rect 246435 397699 246501 397700
rect 245515 397492 245581 397493
rect 245515 397428 245516 397492
rect 245580 397428 245581 397492
rect 245515 397427 245581 397428
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244043 11796 244109 11797
rect 244043 11732 244044 11796
rect 244108 11732 244109 11796
rect 244043 11731 244109 11732
rect 242755 10436 242821 10437
rect 242755 10372 242756 10436
rect 242820 10372 242821 10436
rect 242755 10371 242821 10372
rect 242571 10300 242637 10301
rect 242571 10236 242572 10300
rect 242636 10236 242637 10300
rect 242571 10235 242637 10236
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 -6106 245414 29898
rect 245518 11661 245578 397427
rect 246438 82109 246498 397699
rect 246619 397628 246685 397629
rect 246619 397564 246620 397628
rect 246684 397564 246685 397628
rect 246619 397563 246685 397564
rect 246435 82108 246501 82109
rect 246435 82044 246436 82108
rect 246500 82044 246501 82108
rect 246435 82043 246501 82044
rect 246622 22813 246682 397563
rect 246803 397492 246869 397493
rect 246803 397428 246804 397492
rect 246868 397428 246869 397492
rect 246803 397427 246869 397428
rect 246619 22812 246685 22813
rect 246619 22748 246620 22812
rect 246684 22748 246685 22812
rect 246619 22747 246685 22748
rect 246806 13157 246866 397427
rect 246990 396541 247050 398243
rect 247723 397900 247789 397901
rect 247723 397836 247724 397900
rect 247788 397836 247789 397900
rect 247723 397835 247789 397836
rect 246987 396540 247053 396541
rect 246987 396476 246988 396540
rect 247052 396476 247053 396540
rect 246987 396475 247053 396476
rect 247726 354245 247786 397835
rect 247907 397764 247973 397765
rect 247907 397700 247908 397764
rect 247972 397700 247973 397764
rect 247907 397699 247973 397700
rect 248643 397764 248709 397765
rect 248643 397700 248644 397764
rect 248708 397700 248709 397764
rect 248643 397699 248709 397700
rect 247723 354244 247789 354245
rect 247723 354180 247724 354244
rect 247788 354180 247789 354244
rect 247723 354179 247789 354180
rect 247910 22677 247970 397699
rect 248091 397628 248157 397629
rect 248091 397564 248092 397628
rect 248156 397564 248157 397628
rect 248091 397563 248157 397564
rect 247907 22676 247973 22677
rect 247907 22612 247908 22676
rect 247972 22612 247973 22676
rect 247907 22611 247973 22612
rect 246803 13156 246869 13157
rect 246803 13092 246804 13156
rect 246868 13092 246869 13156
rect 246803 13091 246869 13092
rect 248094 13021 248154 397563
rect 248275 397492 248341 397493
rect 248275 397428 248276 397492
rect 248340 397428 248341 397492
rect 248275 397427 248341 397428
rect 248091 13020 248157 13021
rect 248091 12956 248092 13020
rect 248156 12956 248157 13020
rect 248091 12955 248157 12956
rect 245515 11660 245581 11661
rect 245515 11596 245516 11660
rect 245580 11596 245581 11660
rect 245515 11595 245581 11596
rect 248278 3637 248338 397427
rect 248646 352749 248706 397699
rect 248827 397628 248893 397629
rect 248827 397564 248828 397628
rect 248892 397564 248893 397628
rect 248827 397563 248893 397564
rect 248643 352748 248709 352749
rect 248643 352684 248644 352748
rect 248708 352684 248709 352748
rect 248643 352683 248709 352684
rect 248830 24309 248890 397563
rect 249011 397492 249077 397493
rect 249011 397428 249012 397492
rect 249076 397428 249077 397492
rect 249011 397427 249077 397428
rect 248827 24308 248893 24309
rect 248827 24244 248828 24308
rect 248892 24244 248893 24308
rect 248827 24243 248893 24244
rect 248275 3636 248341 3637
rect 248275 3572 248276 3636
rect 248340 3572 248341 3636
rect 248275 3571 248341 3572
rect 249014 3501 249074 397427
rect 249294 394954 249914 398000
rect 250302 397493 250362 398787
rect 252878 398717 252938 399875
rect 258582 398989 258642 446523
rect 267294 446000 267914 448398
rect 271794 453454 272414 488000
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 264099 445908 264165 445909
rect 264099 445844 264100 445908
rect 264164 445844 264165 445908
rect 264099 445843 264165 445844
rect 262627 445772 262693 445773
rect 262627 445708 262628 445772
rect 262692 445708 262693 445772
rect 262627 445707 262693 445708
rect 262443 444820 262509 444821
rect 262443 444756 262444 444820
rect 262508 444756 262509 444820
rect 262443 444755 262509 444756
rect 261523 444412 261589 444413
rect 261523 444348 261524 444412
rect 261588 444348 261589 444412
rect 261523 444347 261589 444348
rect 260051 444276 260117 444277
rect 260051 444212 260052 444276
rect 260116 444212 260117 444276
rect 260051 444211 260117 444212
rect 260054 401573 260114 444211
rect 261339 443596 261405 443597
rect 261339 443532 261340 443596
rect 261404 443532 261405 443596
rect 261339 443531 261405 443532
rect 260235 441692 260301 441693
rect 260235 441628 260236 441692
rect 260300 441628 260301 441692
rect 260235 441627 260301 441628
rect 260051 401572 260117 401573
rect 260051 401508 260052 401572
rect 260116 401508 260117 401572
rect 260051 401507 260117 401508
rect 258579 398988 258645 398989
rect 258579 398924 258580 398988
rect 258644 398924 258645 398988
rect 258579 398923 258645 398924
rect 260238 398717 260298 441627
rect 252875 398716 252941 398717
rect 252875 398652 252876 398716
rect 252940 398652 252941 398716
rect 252875 398651 252941 398652
rect 260235 398716 260301 398717
rect 260235 398652 260236 398716
rect 260300 398652 260301 398716
rect 260235 398651 260301 398652
rect 253427 398444 253493 398445
rect 253427 398380 253428 398444
rect 253492 398380 253493 398444
rect 253427 398379 253493 398380
rect 250483 397900 250549 397901
rect 250483 397836 250484 397900
rect 250548 397836 250549 397900
rect 250483 397835 250549 397836
rect 251771 397900 251837 397901
rect 251771 397836 251772 397900
rect 251836 397836 251837 397900
rect 251771 397835 251837 397836
rect 250299 397492 250365 397493
rect 250299 397428 250300 397492
rect 250364 397428 250365 397492
rect 250299 397427 250365 397428
rect 250486 395453 250546 397835
rect 250667 397764 250733 397765
rect 250667 397700 250668 397764
rect 250732 397700 250733 397764
rect 250667 397699 250733 397700
rect 250483 395452 250549 395453
rect 250483 395388 250484 395452
rect 250548 395388 250549 395452
rect 250483 395387 250549 395388
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249011 3500 249077 3501
rect 249011 3436 249012 3500
rect 249076 3436 249077 3500
rect 249011 3435 249077 3436
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 -7066 249914 34398
rect 250670 16149 250730 397699
rect 250851 397628 250917 397629
rect 250851 397564 250852 397628
rect 250916 397564 250917 397628
rect 250851 397563 250917 397564
rect 250667 16148 250733 16149
rect 250667 16084 250668 16148
rect 250732 16084 250733 16148
rect 250667 16083 250733 16084
rect 250854 14517 250914 397563
rect 251035 397492 251101 397493
rect 251035 397428 251036 397492
rect 251100 397428 251101 397492
rect 251035 397427 251101 397428
rect 250851 14516 250917 14517
rect 250851 14452 250852 14516
rect 250916 14452 250917 14516
rect 250851 14451 250917 14452
rect 251038 4997 251098 397427
rect 251774 354109 251834 397835
rect 251955 397764 252021 397765
rect 251955 397700 251956 397764
rect 252020 397700 252021 397764
rect 251955 397699 252021 397700
rect 253243 397764 253309 397765
rect 253243 397700 253244 397764
rect 253308 397700 253309 397764
rect 253243 397699 253309 397700
rect 251771 354108 251837 354109
rect 251771 354044 251772 354108
rect 251836 354044 251837 354108
rect 251771 354043 251837 354044
rect 251958 86189 252018 397699
rect 252139 397628 252205 397629
rect 252139 397564 252140 397628
rect 252204 397564 252205 397628
rect 252139 397563 252205 397564
rect 251955 86188 252021 86189
rect 251955 86124 251956 86188
rect 252020 86124 252021 86188
rect 251955 86123 252021 86124
rect 252142 16013 252202 397563
rect 252323 397492 252389 397493
rect 252323 397428 252324 397492
rect 252388 397428 252389 397492
rect 252323 397427 252389 397428
rect 253059 397492 253125 397493
rect 253059 397428 253060 397492
rect 253124 397428 253125 397492
rect 253059 397427 253125 397428
rect 252139 16012 252205 16013
rect 252139 15948 252140 16012
rect 252204 15948 252205 16012
rect 252139 15947 252205 15948
rect 251035 4996 251101 4997
rect 251035 4932 251036 4996
rect 251100 4932 251101 4996
rect 251035 4931 251101 4932
rect 252326 4861 252386 397427
rect 253062 395317 253122 397427
rect 253059 395316 253125 395317
rect 253059 395252 253060 395316
rect 253124 395252 253125 395316
rect 253059 395251 253125 395252
rect 253246 355333 253306 397699
rect 253243 355332 253309 355333
rect 253243 355268 253244 355332
rect 253308 355268 253309 355332
rect 253243 355267 253309 355268
rect 253430 353973 253490 398379
rect 253611 397492 253677 397493
rect 253611 397428 253612 397492
rect 253676 397428 253677 397492
rect 253611 397427 253677 397428
rect 253427 353972 253493 353973
rect 253427 353908 253428 353972
rect 253492 353908 253493 353972
rect 253427 353907 253493 353908
rect 253614 15877 253674 397427
rect 253794 363454 254414 398000
rect 254715 397900 254781 397901
rect 254715 397836 254716 397900
rect 254780 397836 254781 397900
rect 254715 397835 254781 397836
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 254718 352613 254778 397835
rect 254899 397764 254965 397765
rect 254899 397700 254900 397764
rect 254964 397700 254965 397764
rect 254899 397699 254965 397700
rect 254715 352612 254781 352613
rect 254715 352548 254716 352612
rect 254780 352548 254781 352612
rect 254715 352547 254781 352548
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253611 15876 253677 15877
rect 253611 15812 253612 15876
rect 253676 15812 253677 15876
rect 253611 15811 253677 15812
rect 252323 4860 252389 4861
rect 252323 4796 252324 4860
rect 252388 4796 252389 4860
rect 252323 4795 252389 4796
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3454 254414 38898
rect 254902 24173 254962 397699
rect 255083 397628 255149 397629
rect 255083 397564 255084 397628
rect 255148 397564 255149 397628
rect 255083 397563 255149 397564
rect 254899 24172 254965 24173
rect 254899 24108 254900 24172
rect 254964 24108 254965 24172
rect 254899 24107 254965 24108
rect 255086 6221 255146 397563
rect 258294 367954 258914 398000
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 261342 71909 261402 443531
rect 261526 398581 261586 444347
rect 261523 398580 261589 398581
rect 261523 398516 261524 398580
rect 261588 398516 261589 398580
rect 261523 398515 261589 398516
rect 261339 71908 261405 71909
rect 261339 71844 261340 71908
rect 261404 71844 261405 71908
rect 261339 71843 261405 71844
rect 262446 45661 262506 444755
rect 262443 45660 262509 45661
rect 262443 45596 262444 45660
rect 262508 45596 262509 45660
rect 262443 45595 262509 45596
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 255083 6220 255149 6221
rect 255083 6156 255084 6220
rect 255148 6156 255149 6220
rect 255083 6155 255149 6156
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 -1306 258914 7398
rect 262630 3365 262690 445707
rect 264102 398853 264162 445843
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 264099 398852 264165 398853
rect 264099 398788 264100 398852
rect 264164 398788 264165 398852
rect 264099 398787 264165 398788
rect 262794 372454 263414 398000
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262627 3364 262693 3365
rect 262627 3300 262628 3364
rect 262692 3300 262693 3364
rect 262627 3299 262693 3300
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 376954 267914 398000
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 457954 276914 488000
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 462454 281414 488000
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 282134 446453 282194 589867
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 282131 446452 282197 446453
rect 282131 446388 282132 446452
rect 282196 446388 282197 446452
rect 282131 446387 282197 446388
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 691292 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 691292 303914 700398
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 691292 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 691292 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 691292 339914 700398
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 691292 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 691292 371414 695898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 691292 375914 700398
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 300952 687454 301300 687486
rect 300952 687218 301008 687454
rect 301244 687218 301300 687454
rect 300952 687134 301300 687218
rect 300952 686898 301008 687134
rect 301244 686898 301300 687134
rect 300952 686866 301300 686898
rect 389760 687454 390108 687486
rect 389760 687218 389816 687454
rect 390052 687218 390108 687454
rect 389760 687134 390108 687218
rect 389760 686898 389816 687134
rect 390052 686898 390108 687134
rect 389760 686866 390108 686898
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 300272 655954 300620 655986
rect 300272 655718 300328 655954
rect 300564 655718 300620 655954
rect 300272 655634 300620 655718
rect 300272 655398 300328 655634
rect 300564 655398 300620 655634
rect 300272 655366 300620 655398
rect 390440 655954 390788 655986
rect 390440 655718 390496 655954
rect 390732 655718 390788 655954
rect 390440 655634 390788 655718
rect 390440 655398 390496 655634
rect 390732 655398 390788 655634
rect 390440 655366 390788 655398
rect 300952 651454 301300 651486
rect 300952 651218 301008 651454
rect 301244 651218 301300 651454
rect 300952 651134 301300 651218
rect 300952 650898 301008 651134
rect 301244 650898 301300 651134
rect 300952 650866 301300 650898
rect 389760 651454 390108 651486
rect 389760 651218 389816 651454
rect 390052 651218 390108 651454
rect 389760 651134 390108 651218
rect 389760 650898 389816 651134
rect 390052 650898 390108 651134
rect 389760 650866 390108 650898
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 300272 619954 300620 619986
rect 300272 619718 300328 619954
rect 300564 619718 300620 619954
rect 300272 619634 300620 619718
rect 300272 619398 300328 619634
rect 300564 619398 300620 619634
rect 300272 619366 300620 619398
rect 390440 619954 390788 619986
rect 390440 619718 390496 619954
rect 390732 619718 390788 619954
rect 390440 619634 390788 619718
rect 390440 619398 390496 619634
rect 390732 619398 390788 619634
rect 390440 619366 390788 619398
rect 300952 615454 301300 615486
rect 300952 615218 301008 615454
rect 301244 615218 301300 615454
rect 300952 615134 301300 615218
rect 300952 614898 301008 615134
rect 301244 614898 301300 615134
rect 300952 614866 301300 614898
rect 389760 615454 390108 615486
rect 389760 615218 389816 615454
rect 390052 615218 390108 615454
rect 389760 615134 390108 615218
rect 389760 614898 389816 615134
rect 390052 614898 390108 615134
rect 389760 614866 390108 614898
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 312928 599450 312988 600100
rect 312862 599390 312988 599450
rect 314288 599450 314348 600100
rect 315376 599450 315436 600100
rect 317688 599586 317748 600100
rect 314288 599390 314394 599450
rect 312862 596597 312922 599390
rect 314334 597277 314394 599390
rect 315254 599390 315436 599450
rect 317646 599526 317748 599586
rect 318912 599586 318972 600100
rect 320000 599586 320060 600100
rect 321088 599586 321148 600100
rect 322312 599586 322372 600100
rect 323400 599586 323460 600100
rect 318912 599526 318994 599586
rect 320000 599526 320098 599586
rect 321088 599526 321202 599586
rect 314331 597276 314397 597277
rect 314331 597212 314332 597276
rect 314396 597212 314397 597276
rect 314331 597211 314397 597212
rect 315254 596869 315314 599390
rect 317646 597549 317706 599526
rect 317643 597548 317709 597549
rect 317643 597484 317644 597548
rect 317708 597484 317709 597548
rect 317643 597483 317709 597484
rect 318934 597413 318994 599526
rect 320038 597549 320098 599526
rect 321142 597549 321202 599526
rect 322246 599526 322372 599586
rect 323350 599526 323460 599586
rect 324760 599586 324820 600100
rect 325304 599586 325364 600100
rect 324760 599526 324882 599586
rect 322246 597549 322306 599526
rect 323350 597549 323410 599526
rect 320035 597548 320101 597549
rect 320035 597484 320036 597548
rect 320100 597484 320101 597548
rect 320035 597483 320101 597484
rect 321139 597548 321205 597549
rect 321139 597484 321140 597548
rect 321204 597484 321205 597548
rect 321139 597483 321205 597484
rect 322243 597548 322309 597549
rect 322243 597484 322244 597548
rect 322308 597484 322309 597548
rect 322243 597483 322309 597484
rect 323347 597548 323413 597549
rect 323347 597484 323348 597548
rect 323412 597484 323413 597548
rect 323347 597483 323413 597484
rect 324822 597413 324882 599526
rect 325190 599526 325364 599586
rect 325712 599586 325772 600100
rect 330472 599586 330532 600100
rect 325712 599526 325802 599586
rect 330472 599526 330586 599586
rect 325190 597549 325250 599526
rect 325742 597549 325802 599526
rect 330526 597549 330586 599526
rect 335504 599450 335564 600100
rect 340536 599450 340596 600100
rect 335126 599390 335564 599450
rect 340462 599390 340596 599450
rect 345568 599450 345628 600100
rect 350464 599450 350524 600100
rect 355496 599450 355556 600100
rect 360528 599450 360588 600100
rect 345568 599390 345674 599450
rect 325187 597548 325253 597549
rect 325187 597484 325188 597548
rect 325252 597484 325253 597548
rect 325187 597483 325253 597484
rect 325739 597548 325805 597549
rect 325739 597484 325740 597548
rect 325804 597484 325805 597548
rect 325739 597483 325805 597484
rect 330523 597548 330589 597549
rect 330523 597484 330524 597548
rect 330588 597484 330589 597548
rect 330523 597483 330589 597484
rect 335126 597413 335186 599390
rect 318931 597412 318997 597413
rect 318931 597348 318932 597412
rect 318996 597348 318997 597412
rect 318931 597347 318997 597348
rect 324819 597412 324885 597413
rect 324819 597348 324820 597412
rect 324884 597348 324885 597412
rect 324819 597347 324885 597348
rect 335123 597412 335189 597413
rect 335123 597348 335124 597412
rect 335188 597348 335189 597412
rect 335123 597347 335189 597348
rect 340462 597005 340522 599390
rect 345614 597549 345674 599390
rect 350398 599390 350524 599450
rect 354446 599390 355556 599450
rect 360518 599390 360588 599450
rect 345611 597548 345677 597549
rect 345611 597484 345612 597548
rect 345676 597484 345677 597548
rect 345611 597483 345677 597484
rect 350398 597141 350458 599390
rect 350395 597140 350461 597141
rect 350395 597076 350396 597140
rect 350460 597076 350461 597140
rect 350395 597075 350461 597076
rect 340459 597004 340525 597005
rect 340459 596940 340460 597004
rect 340524 596940 340525 597004
rect 340459 596939 340525 596940
rect 315251 596868 315317 596869
rect 315251 596804 315252 596868
rect 315316 596804 315317 596868
rect 315251 596803 315317 596804
rect 312859 596596 312925 596597
rect 312859 596532 312860 596596
rect 312924 596532 312925 596596
rect 312859 596531 312925 596532
rect 354446 596325 354506 599390
rect 360518 597549 360578 599390
rect 360515 597548 360581 597549
rect 360515 597484 360516 597548
rect 360580 597484 360581 597548
rect 360515 597483 360581 597484
rect 354443 596324 354509 596325
rect 354443 596260 354444 596324
rect 354508 596260 354509 596324
rect 354443 596259 354509 596260
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 300272 547954 300620 547986
rect 300272 547718 300328 547954
rect 300564 547718 300620 547954
rect 300272 547634 300620 547718
rect 300272 547398 300328 547634
rect 300564 547398 300620 547634
rect 300272 547366 300620 547398
rect 390440 547954 390788 547986
rect 390440 547718 390496 547954
rect 390732 547718 390788 547954
rect 390440 547634 390788 547718
rect 390440 547398 390496 547634
rect 390732 547398 390788 547634
rect 390440 547366 390788 547398
rect 300952 543454 301300 543486
rect 300952 543218 301008 543454
rect 301244 543218 301300 543454
rect 300952 543134 301300 543218
rect 300952 542898 301008 543134
rect 301244 542898 301300 543134
rect 300952 542866 301300 542898
rect 389760 543454 390108 543486
rect 389760 543218 389816 543454
rect 390052 543218 390108 543454
rect 389760 543134 390108 543218
rect 389760 542898 389816 543134
rect 390052 542898 390108 543134
rect 389760 542866 390108 542898
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 300272 511954 300620 511986
rect 300272 511718 300328 511954
rect 300564 511718 300620 511954
rect 300272 511634 300620 511718
rect 300272 511398 300328 511634
rect 300564 511398 300620 511634
rect 300272 511366 300620 511398
rect 390440 511954 390788 511986
rect 390440 511718 390496 511954
rect 390732 511718 390788 511954
rect 390440 511634 390788 511718
rect 390440 511398 390496 511634
rect 390732 511398 390788 511634
rect 390440 511366 390788 511398
rect 300952 507454 301300 507486
rect 300952 507218 301008 507454
rect 301244 507218 301300 507454
rect 300952 507134 301300 507218
rect 300952 506898 301008 507134
rect 301244 506898 301300 507134
rect 300952 506866 301300 506898
rect 389760 507454 390108 507486
rect 389760 507218 389816 507454
rect 390052 507218 390108 507454
rect 389760 507134 390108 507218
rect 389760 506898 389816 507134
rect 390052 506898 390108 507134
rect 389760 506866 390108 506898
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 312928 489930 312988 490106
rect 314288 489930 314348 490106
rect 315376 489930 315436 490106
rect 317688 489930 317748 490106
rect 312928 489870 313106 489930
rect 314288 489870 314394 489930
rect 315376 489870 315498 489930
rect 313046 487933 313106 489870
rect 314334 488477 314394 489870
rect 315438 488477 315498 489870
rect 317646 489870 317748 489930
rect 318912 489930 318972 490106
rect 320000 489930 320060 490106
rect 321088 489930 321148 490106
rect 322312 489930 322372 490106
rect 323400 489930 323460 490106
rect 324760 489930 324820 490106
rect 325304 489930 325364 490106
rect 318912 489870 318994 489930
rect 320000 489870 320098 489930
rect 321088 489870 321202 489930
rect 314331 488476 314397 488477
rect 314331 488412 314332 488476
rect 314396 488412 314397 488476
rect 314331 488411 314397 488412
rect 315435 488476 315501 488477
rect 315435 488412 315436 488476
rect 315500 488412 315501 488476
rect 315435 488411 315501 488412
rect 313043 487932 313109 487933
rect 313043 487868 313044 487932
rect 313108 487868 313109 487932
rect 313043 487867 313109 487868
rect 317646 487253 317706 489870
rect 318934 487253 318994 489870
rect 320038 487525 320098 489870
rect 320035 487524 320101 487525
rect 320035 487460 320036 487524
rect 320100 487460 320101 487524
rect 320035 487459 320101 487460
rect 321142 487253 321202 489870
rect 322246 489870 322372 489930
rect 323350 489870 323460 489930
rect 324638 489870 324820 489930
rect 325190 489870 325364 489930
rect 325712 489930 325772 490106
rect 330472 489930 330532 490106
rect 335504 489930 335564 490106
rect 340536 489930 340596 490106
rect 325712 489870 325802 489930
rect 330472 489870 330586 489930
rect 322246 487389 322306 489870
rect 323350 487525 323410 489870
rect 324638 487933 324698 489870
rect 324635 487932 324701 487933
rect 324635 487868 324636 487932
rect 324700 487868 324701 487932
rect 324635 487867 324701 487868
rect 323347 487524 323413 487525
rect 323347 487460 323348 487524
rect 323412 487460 323413 487524
rect 323347 487459 323413 487460
rect 322243 487388 322309 487389
rect 322243 487324 322244 487388
rect 322308 487324 322309 487388
rect 322243 487323 322309 487324
rect 325190 487253 325250 489870
rect 325742 487797 325802 489870
rect 325739 487796 325805 487797
rect 325739 487732 325740 487796
rect 325804 487732 325805 487796
rect 325739 487731 325805 487732
rect 330526 487253 330586 489870
rect 335494 489870 335564 489930
rect 340462 489870 340596 489930
rect 345568 489930 345628 490106
rect 350464 489930 350524 490106
rect 345568 489870 345674 489930
rect 335494 487253 335554 489870
rect 340462 487253 340522 489870
rect 345614 487253 345674 489870
rect 350398 489870 350524 489930
rect 355496 489930 355556 490106
rect 360528 489930 360588 490106
rect 355496 489870 355610 489930
rect 350398 487253 350458 489870
rect 355550 487253 355610 489870
rect 360518 489870 360588 489930
rect 360518 487253 360578 489870
rect 317643 487252 317709 487253
rect 317643 487188 317644 487252
rect 317708 487188 317709 487252
rect 317643 487187 317709 487188
rect 318931 487252 318997 487253
rect 318931 487188 318932 487252
rect 318996 487188 318997 487252
rect 318931 487187 318997 487188
rect 321139 487252 321205 487253
rect 321139 487188 321140 487252
rect 321204 487188 321205 487252
rect 321139 487187 321205 487188
rect 325187 487252 325253 487253
rect 325187 487188 325188 487252
rect 325252 487188 325253 487252
rect 325187 487187 325253 487188
rect 330523 487252 330589 487253
rect 330523 487188 330524 487252
rect 330588 487188 330589 487252
rect 330523 487187 330589 487188
rect 335491 487252 335557 487253
rect 335491 487188 335492 487252
rect 335556 487188 335557 487252
rect 335491 487187 335557 487188
rect 340459 487252 340525 487253
rect 340459 487188 340460 487252
rect 340524 487188 340525 487252
rect 340459 487187 340525 487188
rect 345611 487252 345677 487253
rect 345611 487188 345612 487252
rect 345676 487188 345677 487252
rect 345611 487187 345677 487188
rect 350395 487252 350461 487253
rect 350395 487188 350396 487252
rect 350460 487188 350461 487252
rect 350395 487187 350461 487188
rect 355547 487252 355613 487253
rect 355547 487188 355548 487252
rect 355612 487188 355613 487252
rect 355547 487187 355613 487188
rect 360515 487252 360581 487253
rect 360515 487188 360516 487252
rect 360580 487188 360581 487252
rect 360515 487187 360581 487188
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 293171 448764 293237 448765
rect 293171 448700 293172 448764
rect 293236 448700 293237 448764
rect 293171 448699 293237 448700
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 293174 397901 293234 448699
rect 294294 439954 294914 475398
rect 388794 462454 389414 488000
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 382227 454340 382293 454341
rect 382227 454276 382228 454340
rect 382292 454276 382293 454340
rect 382227 454275 382293 454276
rect 298507 446180 298573 446181
rect 298507 446116 298508 446180
rect 298572 446116 298573 446180
rect 298507 446115 298573 446116
rect 295931 442236 295997 442237
rect 295931 442172 295932 442236
rect 295996 442172 295997 442236
rect 295931 442171 295997 442172
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 293171 397900 293237 397901
rect 293171 397836 293172 397900
rect 293236 397836 293237 397900
rect 293171 397835 293237 397836
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 295934 19413 295994 442171
rect 295931 19412 295997 19413
rect 295931 19348 295932 19412
rect 295996 19348 295997 19412
rect 295931 19347 295997 19348
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 298510 5677 298570 446115
rect 319568 439954 319888 439986
rect 319568 439718 319610 439954
rect 319846 439718 319888 439954
rect 319568 439634 319888 439718
rect 319568 439398 319610 439634
rect 319846 439398 319888 439634
rect 319568 439366 319888 439398
rect 350288 439954 350608 439986
rect 350288 439718 350330 439954
rect 350566 439718 350608 439954
rect 350288 439634 350608 439718
rect 350288 439398 350330 439634
rect 350566 439398 350608 439634
rect 350288 439366 350608 439398
rect 381008 439954 381328 439986
rect 381008 439718 381050 439954
rect 381286 439718 381328 439954
rect 381008 439634 381328 439718
rect 381008 439398 381050 439634
rect 381286 439398 381328 439634
rect 381008 439366 381328 439398
rect 304208 435454 304528 435486
rect 304208 435218 304250 435454
rect 304486 435218 304528 435454
rect 304208 435134 304528 435218
rect 304208 434898 304250 435134
rect 304486 434898 304528 435134
rect 304208 434866 304528 434898
rect 334928 435454 335248 435486
rect 334928 435218 334970 435454
rect 335206 435218 335248 435454
rect 334928 435134 335248 435218
rect 334928 434898 334970 435134
rect 335206 434898 335248 435134
rect 334928 434866 335248 434898
rect 365648 435454 365968 435486
rect 365648 435218 365690 435454
rect 365926 435218 365968 435454
rect 365648 435134 365968 435218
rect 365648 434898 365690 435134
rect 365926 434898 365968 435134
rect 365648 434866 365968 434898
rect 382230 422310 382290 454275
rect 382411 454204 382477 454205
rect 382411 454140 382412 454204
rect 382476 454140 382477 454204
rect 382411 454139 382477 454140
rect 382414 441630 382474 454139
rect 382414 441570 383394 441630
rect 383334 425781 383394 441570
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 383331 425780 383397 425781
rect 383331 425716 383332 425780
rect 383396 425716 383397 425780
rect 383331 425715 383397 425716
rect 382230 422250 383394 422310
rect 383334 412589 383394 422250
rect 383331 412588 383397 412589
rect 383331 412524 383332 412588
rect 383396 412524 383397 412588
rect 383331 412523 383397 412524
rect 319568 403954 319888 403986
rect 319568 403718 319610 403954
rect 319846 403718 319888 403954
rect 319568 403634 319888 403718
rect 319568 403398 319610 403634
rect 319846 403398 319888 403634
rect 319568 403366 319888 403398
rect 350288 403954 350608 403986
rect 350288 403718 350330 403954
rect 350566 403718 350608 403954
rect 350288 403634 350608 403718
rect 350288 403398 350330 403634
rect 350566 403398 350608 403634
rect 350288 403366 350608 403398
rect 381008 403954 381328 403986
rect 381008 403718 381050 403954
rect 381286 403718 381328 403954
rect 381008 403634 381328 403718
rect 381008 403398 381050 403634
rect 381286 403398 381328 403634
rect 381008 403366 381328 403398
rect 383331 402932 383397 402933
rect 383331 402868 383332 402932
rect 383396 402868 383397 402932
rect 383331 402867 383397 402868
rect 383334 401573 383394 402867
rect 383331 401572 383397 401573
rect 383331 401508 383332 401572
rect 383396 401508 383397 401572
rect 383331 401507 383397 401508
rect 298794 372454 299414 398000
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 5676 298573 5677
rect 298507 5612 298508 5676
rect 298572 5612 298573 5676
rect 298507 5611 298573 5612
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 376954 303914 398000
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 381454 308414 398000
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 385954 312914 398000
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 390454 317414 398000
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 394954 321914 398000
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 367954 330914 398000
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 372454 335414 398000
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 376954 339914 398000
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 385954 348914 398000
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 390454 353414 398000
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 394954 357914 398000
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 363454 362414 398000
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 367954 366914 398000
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 372454 371414 398000
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 376954 375914 398000
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 381454 380414 398000
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 385954 384914 398000
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 691292 411914 700398
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 691292 438914 691398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 691292 443414 695898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 691292 447914 700398
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 691292 474914 691398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 691292 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 691292 483914 700398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 410952 687454 411300 687486
rect 410952 687218 411008 687454
rect 411244 687218 411300 687454
rect 410952 687134 411300 687218
rect 410952 686898 411008 687134
rect 411244 686898 411300 687134
rect 410952 686866 411300 686898
rect 499760 687454 500108 687486
rect 499760 687218 499816 687454
rect 500052 687218 500108 687454
rect 499760 687134 500108 687218
rect 499760 686898 499816 687134
rect 500052 686898 500108 687134
rect 499760 686866 500108 686898
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 410272 655954 410620 655986
rect 410272 655718 410328 655954
rect 410564 655718 410620 655954
rect 410272 655634 410620 655718
rect 410272 655398 410328 655634
rect 410564 655398 410620 655634
rect 410272 655366 410620 655398
rect 500440 655954 500788 655986
rect 500440 655718 500496 655954
rect 500732 655718 500788 655954
rect 500440 655634 500788 655718
rect 500440 655398 500496 655634
rect 500732 655398 500788 655634
rect 500440 655366 500788 655398
rect 410952 651454 411300 651486
rect 410952 651218 411008 651454
rect 411244 651218 411300 651454
rect 410952 651134 411300 651218
rect 410952 650898 411008 651134
rect 411244 650898 411300 651134
rect 410952 650866 411300 650898
rect 499760 651454 500108 651486
rect 499760 651218 499816 651454
rect 500052 651218 500108 651454
rect 499760 651134 500108 651218
rect 499760 650898 499816 651134
rect 500052 650898 500108 651134
rect 499760 650866 500108 650898
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 410272 619954 410620 619986
rect 410272 619718 410328 619954
rect 410564 619718 410620 619954
rect 410272 619634 410620 619718
rect 410272 619398 410328 619634
rect 410564 619398 410620 619634
rect 410272 619366 410620 619398
rect 500440 619954 500788 619986
rect 500440 619718 500496 619954
rect 500732 619718 500788 619954
rect 500440 619634 500788 619718
rect 500440 619398 500496 619634
rect 500732 619398 500788 619634
rect 500440 619366 500788 619398
rect 410952 615454 411300 615486
rect 410952 615218 411008 615454
rect 411244 615218 411300 615454
rect 410952 615134 411300 615218
rect 410952 614898 411008 615134
rect 411244 614898 411300 615134
rect 410952 614866 411300 614898
rect 499760 615454 500108 615486
rect 499760 615218 499816 615454
rect 500052 615218 500108 615454
rect 499760 615134 500108 615218
rect 499760 614898 499816 615134
rect 500052 614898 500108 615134
rect 499760 614866 500108 614898
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 422928 599450 422988 600100
rect 424288 599450 424348 600100
rect 425376 599450 425436 600100
rect 427688 599450 427748 600100
rect 422894 599390 422988 599450
rect 424182 599390 424348 599450
rect 425286 599390 425436 599450
rect 427678 599390 427748 599450
rect 428912 599450 428972 600100
rect 430000 599450 430060 600100
rect 431088 599450 431148 600100
rect 432312 599450 432372 600100
rect 433400 599450 433460 600100
rect 434760 599450 434820 600100
rect 435304 599450 435364 600100
rect 435712 599450 435772 600100
rect 440472 599450 440532 600100
rect 428912 599390 429026 599450
rect 422894 597277 422954 599390
rect 422891 597276 422957 597277
rect 422891 597212 422892 597276
rect 422956 597212 422957 597276
rect 422891 597211 422957 597212
rect 424182 597005 424242 599390
rect 424179 597004 424245 597005
rect 424179 596940 424180 597004
rect 424244 596940 424245 597004
rect 424179 596939 424245 596940
rect 425286 596461 425346 599390
rect 427678 597277 427738 599390
rect 428966 597413 429026 599390
rect 429886 599390 430060 599450
rect 430990 599390 431148 599450
rect 431726 599390 432372 599450
rect 433382 599390 433460 599450
rect 434670 599390 434820 599450
rect 435222 599390 435364 599450
rect 435590 599390 435772 599450
rect 440374 599390 440532 599450
rect 445504 599450 445564 600100
rect 450536 599450 450596 600100
rect 455568 599450 455628 600100
rect 460464 599450 460524 600100
rect 465496 599450 465556 600100
rect 470528 599450 470588 600100
rect 445504 599390 445586 599450
rect 428963 597412 429029 597413
rect 428963 597348 428964 597412
rect 429028 597348 429029 597412
rect 428963 597347 429029 597348
rect 427675 597276 427741 597277
rect 427675 597212 427676 597276
rect 427740 597212 427741 597276
rect 427675 597211 427741 597212
rect 429886 597005 429946 599390
rect 430990 597413 431050 599390
rect 430987 597412 431053 597413
rect 430987 597348 430988 597412
rect 431052 597348 431053 597412
rect 430987 597347 431053 597348
rect 431726 597005 431786 599390
rect 433382 597141 433442 599390
rect 434670 597141 434730 599390
rect 433379 597140 433445 597141
rect 433379 597076 433380 597140
rect 433444 597076 433445 597140
rect 433379 597075 433445 597076
rect 434667 597140 434733 597141
rect 434667 597076 434668 597140
rect 434732 597076 434733 597140
rect 434667 597075 434733 597076
rect 429883 597004 429949 597005
rect 429883 596940 429884 597004
rect 429948 596940 429949 597004
rect 429883 596939 429949 596940
rect 431723 597004 431789 597005
rect 431723 596940 431724 597004
rect 431788 596940 431789 597004
rect 431723 596939 431789 596940
rect 435222 596733 435282 599390
rect 435590 597413 435650 599390
rect 440374 597549 440434 599390
rect 440371 597548 440437 597549
rect 440371 597484 440372 597548
rect 440436 597484 440437 597548
rect 440371 597483 440437 597484
rect 435587 597412 435653 597413
rect 435587 597348 435588 597412
rect 435652 597348 435653 597412
rect 435587 597347 435653 597348
rect 445526 596733 445586 599390
rect 450494 599390 450596 599450
rect 455462 599390 455628 599450
rect 460430 599390 460524 599450
rect 465398 599390 465556 599450
rect 470366 599390 470588 599450
rect 450494 597549 450554 599390
rect 450491 597548 450557 597549
rect 450491 597484 450492 597548
rect 450556 597484 450557 597548
rect 450491 597483 450557 597484
rect 435219 596732 435285 596733
rect 435219 596668 435220 596732
rect 435284 596668 435285 596732
rect 435219 596667 435285 596668
rect 445523 596732 445589 596733
rect 445523 596668 445524 596732
rect 445588 596668 445589 596732
rect 445523 596667 445589 596668
rect 425283 596460 425349 596461
rect 425283 596396 425284 596460
rect 425348 596396 425349 596460
rect 425283 596395 425349 596396
rect 455462 596325 455522 599390
rect 460430 597549 460490 599390
rect 460427 597548 460493 597549
rect 460427 597484 460428 597548
rect 460492 597484 460493 597548
rect 460427 597483 460493 597484
rect 465398 596869 465458 599390
rect 465395 596868 465461 596869
rect 465395 596804 465396 596868
rect 465460 596804 465461 596868
rect 465395 596803 465461 596804
rect 470366 596325 470426 599390
rect 455459 596324 455525 596325
rect 455459 596260 455460 596324
rect 455524 596260 455525 596324
rect 455459 596259 455525 596260
rect 470363 596324 470429 596325
rect 470363 596260 470364 596324
rect 470428 596260 470429 596324
rect 470363 596259 470429 596260
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 410272 547954 410620 547986
rect 410272 547718 410328 547954
rect 410564 547718 410620 547954
rect 410272 547634 410620 547718
rect 410272 547398 410328 547634
rect 410564 547398 410620 547634
rect 410272 547366 410620 547398
rect 500440 547954 500788 547986
rect 500440 547718 500496 547954
rect 500732 547718 500788 547954
rect 500440 547634 500788 547718
rect 500440 547398 500496 547634
rect 500732 547398 500788 547634
rect 500440 547366 500788 547398
rect 410952 543454 411300 543486
rect 410952 543218 411008 543454
rect 411244 543218 411300 543454
rect 410952 543134 411300 543218
rect 410952 542898 411008 543134
rect 411244 542898 411300 543134
rect 410952 542866 411300 542898
rect 499760 543454 500108 543486
rect 499760 543218 499816 543454
rect 500052 543218 500108 543454
rect 499760 543134 500108 543218
rect 499760 542898 499816 543134
rect 500052 542898 500108 543134
rect 499760 542866 500108 542898
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 407803 526692 407869 526693
rect 407803 526628 407804 526692
rect 407868 526628 407869 526692
rect 407803 526627 407869 526628
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 407806 488069 407866 526627
rect 408171 523700 408237 523701
rect 408171 523636 408172 523700
rect 408236 523636 408237 523700
rect 408171 523635 408237 523636
rect 408174 489837 408234 523635
rect 410272 511954 410620 511986
rect 410272 511718 410328 511954
rect 410564 511718 410620 511954
rect 410272 511634 410620 511718
rect 410272 511398 410328 511634
rect 410564 511398 410620 511634
rect 410272 511366 410620 511398
rect 500440 511954 500788 511986
rect 500440 511718 500496 511954
rect 500732 511718 500788 511954
rect 500440 511634 500788 511718
rect 500440 511398 500496 511634
rect 500732 511398 500788 511634
rect 500440 511366 500788 511398
rect 410952 507454 411300 507486
rect 410952 507218 411008 507454
rect 411244 507218 411300 507454
rect 410952 507134 411300 507218
rect 410952 506898 411008 507134
rect 411244 506898 411300 507134
rect 410952 506866 411300 506898
rect 499760 507454 500108 507486
rect 499760 507218 499816 507454
rect 500052 507218 500108 507454
rect 499760 507134 500108 507218
rect 499760 506898 499816 507134
rect 500052 506898 500108 507134
rect 499760 506866 500108 506898
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 422928 489930 422988 490106
rect 424288 489930 424348 490106
rect 425376 489930 425436 490106
rect 427688 489930 427748 490106
rect 422894 489870 422988 489930
rect 424182 489870 424348 489930
rect 425286 489870 425436 489930
rect 427678 489870 427748 489930
rect 428912 489930 428972 490106
rect 430000 489930 430060 490106
rect 431088 489930 431148 490106
rect 432312 489930 432372 490106
rect 433400 489930 433460 490106
rect 428912 489870 429026 489930
rect 408171 489836 408237 489837
rect 408171 489772 408172 489836
rect 408236 489772 408237 489836
rect 408171 489771 408237 489772
rect 422894 488477 422954 489870
rect 424182 488477 424242 489870
rect 425286 488477 425346 489870
rect 422891 488476 422957 488477
rect 422891 488412 422892 488476
rect 422956 488412 422957 488476
rect 422891 488411 422957 488412
rect 424179 488476 424245 488477
rect 424179 488412 424180 488476
rect 424244 488412 424245 488476
rect 424179 488411 424245 488412
rect 425283 488476 425349 488477
rect 425283 488412 425284 488476
rect 425348 488412 425349 488476
rect 425283 488411 425349 488412
rect 407803 488068 407869 488069
rect 407803 488004 407804 488068
rect 407868 488004 407869 488068
rect 407803 488003 407869 488004
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 484954 411914 488000
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 453454 416414 488000
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 457954 420914 488000
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 462454 425414 488000
rect 427678 487661 427738 489870
rect 428966 487661 429026 489870
rect 429886 489870 430060 489930
rect 430990 489870 431148 489930
rect 432278 489870 432372 489930
rect 433382 489870 433460 489930
rect 434760 489930 434820 490106
rect 435304 489930 435364 490106
rect 435712 489930 435772 490106
rect 440472 489930 440532 490106
rect 434760 489870 434914 489930
rect 429886 488205 429946 489870
rect 429883 488204 429949 488205
rect 429883 488140 429884 488204
rect 429948 488140 429949 488204
rect 429883 488139 429949 488140
rect 427675 487660 427741 487661
rect 427675 487596 427676 487660
rect 427740 487596 427741 487660
rect 427675 487595 427741 487596
rect 428963 487660 429029 487661
rect 428963 487596 428964 487660
rect 429028 487596 429029 487660
rect 428963 487595 429029 487596
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 466954 429914 488000
rect 430990 487797 431050 489870
rect 430987 487796 431053 487797
rect 430987 487732 430988 487796
rect 431052 487732 431053 487796
rect 430987 487731 431053 487732
rect 432278 487389 432338 489870
rect 433382 487525 433442 489870
rect 433379 487524 433445 487525
rect 433379 487460 433380 487524
rect 433444 487460 433445 487524
rect 433379 487459 433445 487460
rect 432275 487388 432341 487389
rect 432275 487324 432276 487388
rect 432340 487324 432341 487388
rect 432275 487323 432341 487324
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 471454 434414 488000
rect 434854 487389 434914 489870
rect 435222 489870 435364 489930
rect 435590 489870 435772 489930
rect 440374 489870 440532 489930
rect 445504 489930 445564 490106
rect 450536 489930 450596 490106
rect 455568 489930 455628 490106
rect 460464 489930 460524 490106
rect 465496 489930 465556 490106
rect 445504 489870 445586 489930
rect 434851 487388 434917 487389
rect 434851 487324 434852 487388
rect 434916 487324 434917 487388
rect 434851 487323 434917 487324
rect 435222 487253 435282 489870
rect 435590 488205 435650 489870
rect 435587 488204 435653 488205
rect 435587 488140 435588 488204
rect 435652 488140 435653 488204
rect 435587 488139 435653 488140
rect 435219 487252 435285 487253
rect 435219 487188 435220 487252
rect 435284 487188 435285 487252
rect 435219 487187 435285 487188
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 475954 438914 488000
rect 440374 487253 440434 489870
rect 440371 487252 440437 487253
rect 440371 487188 440372 487252
rect 440436 487188 440437 487252
rect 440371 487187 440437 487188
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 480454 443414 488000
rect 445526 487253 445586 489870
rect 450494 489870 450596 489930
rect 455462 489870 455628 489930
rect 460430 489870 460524 489930
rect 465398 489870 465556 489930
rect 470528 489930 470588 490106
rect 470528 489870 470794 489930
rect 445523 487252 445589 487253
rect 445523 487188 445524 487252
rect 445588 487188 445589 487252
rect 445523 487187 445589 487188
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 484954 447914 488000
rect 450494 487253 450554 489870
rect 450491 487252 450557 487253
rect 450491 487188 450492 487252
rect 450556 487188 450557 487252
rect 450491 487187 450557 487188
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 453454 452414 488000
rect 455462 487253 455522 489870
rect 455459 487252 455525 487253
rect 455459 487188 455460 487252
rect 455524 487188 455525 487252
rect 455459 487187 455525 487188
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 457954 456914 488000
rect 460430 487253 460490 489870
rect 465398 488341 465458 489870
rect 465395 488340 465461 488341
rect 465395 488276 465396 488340
rect 465460 488276 465461 488340
rect 465395 488275 465461 488276
rect 460427 487252 460493 487253
rect 460427 487188 460428 487252
rect 460492 487188 460493 487252
rect 460427 487187 460493 487188
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 462454 461414 488000
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 466954 465914 488000
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 471454 470414 488000
rect 470734 487253 470794 489870
rect 470731 487252 470797 487253
rect 470731 487188 470732 487252
rect 470796 487188 470797 487252
rect 470731 487187 470797 487188
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 475954 474914 488000
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 480454 479414 488000
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 484954 483914 488000
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 453454 488414 488000
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 457954 492914 488000
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 462454 497414 488000
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 466954 501914 488000
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 81008 687218 81244 687454
rect 81008 686898 81244 687134
rect 169816 687218 170052 687454
rect 169816 686898 170052 687134
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 80328 655718 80564 655954
rect 80328 655398 80564 655634
rect 170496 655718 170732 655954
rect 170496 655398 170732 655634
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 81008 651218 81244 651454
rect 81008 650898 81244 651134
rect 169816 651218 170052 651454
rect 169816 650898 170052 651134
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 80328 619718 80564 619954
rect 80328 619398 80564 619634
rect 170496 619718 170732 619954
rect 170496 619398 170732 619634
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 81008 615218 81244 615454
rect 81008 614898 81244 615134
rect 169816 615218 170052 615454
rect 169816 614898 170052 615134
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 80328 547718 80564 547954
rect 80328 547398 80564 547634
rect 170496 547718 170732 547954
rect 170496 547398 170732 547634
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 81008 543218 81244 543454
rect 81008 542898 81244 543134
rect 169816 543218 170052 543454
rect 169816 542898 170052 543134
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 80328 511718 80564 511954
rect 80328 511398 80564 511634
rect 170496 511718 170732 511954
rect 170496 511398 170732 511634
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 81008 507218 81244 507454
rect 81008 506898 81244 507134
rect 169816 507218 170052 507454
rect 169816 506898 170052 507134
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 191008 687218 191244 687454
rect 191008 686898 191244 687134
rect 279816 687218 280052 687454
rect 279816 686898 280052 687134
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 190328 655718 190564 655954
rect 190328 655398 190564 655634
rect 280496 655718 280732 655954
rect 280496 655398 280732 655634
rect 191008 651218 191244 651454
rect 191008 650898 191244 651134
rect 279816 651218 280052 651454
rect 279816 650898 280052 651134
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190328 619718 190564 619954
rect 190328 619398 190564 619634
rect 280496 619718 280732 619954
rect 280496 619398 280732 619634
rect 191008 615218 191244 615454
rect 191008 614898 191244 615134
rect 279816 615218 280052 615454
rect 279816 614898 280052 615134
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 190328 547718 190564 547954
rect 190328 547398 190564 547634
rect 280496 547718 280732 547954
rect 280496 547398 280732 547634
rect 191008 543218 191244 543454
rect 191008 542898 191244 543134
rect 279816 543218 280052 543454
rect 279816 542898 280052 543134
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 190328 511718 190564 511954
rect 190328 511398 190564 511634
rect 280496 511718 280732 511954
rect 280496 511398 280732 511634
rect 191008 507218 191244 507454
rect 191008 506898 191244 507134
rect 279816 507218 280052 507454
rect 279816 506898 280052 507134
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 219610 439718 219846 439954
rect 219610 439398 219846 439634
rect 250330 439718 250566 439954
rect 250330 439398 250566 439634
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 219610 403718 219846 403954
rect 219610 403398 219846 403634
rect 250330 403718 250566 403954
rect 250330 403398 250566 403634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 301008 687218 301244 687454
rect 301008 686898 301244 687134
rect 389816 687218 390052 687454
rect 389816 686898 390052 687134
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 300328 655718 300564 655954
rect 300328 655398 300564 655634
rect 390496 655718 390732 655954
rect 390496 655398 390732 655634
rect 301008 651218 301244 651454
rect 301008 650898 301244 651134
rect 389816 651218 390052 651454
rect 389816 650898 390052 651134
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 300328 619718 300564 619954
rect 300328 619398 300564 619634
rect 390496 619718 390732 619954
rect 390496 619398 390732 619634
rect 301008 615218 301244 615454
rect 301008 614898 301244 615134
rect 389816 615218 390052 615454
rect 389816 614898 390052 615134
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 300328 547718 300564 547954
rect 300328 547398 300564 547634
rect 390496 547718 390732 547954
rect 390496 547398 390732 547634
rect 301008 543218 301244 543454
rect 301008 542898 301244 543134
rect 389816 543218 390052 543454
rect 389816 542898 390052 543134
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 300328 511718 300564 511954
rect 300328 511398 300564 511634
rect 390496 511718 390732 511954
rect 390496 511398 390732 511634
rect 301008 507218 301244 507454
rect 301008 506898 301244 507134
rect 389816 507218 390052 507454
rect 389816 506898 390052 507134
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 319610 439718 319846 439954
rect 319610 439398 319846 439634
rect 350330 439718 350566 439954
rect 350330 439398 350566 439634
rect 381050 439718 381286 439954
rect 381050 439398 381286 439634
rect 304250 435218 304486 435454
rect 304250 434898 304486 435134
rect 334970 435218 335206 435454
rect 334970 434898 335206 435134
rect 365690 435218 365926 435454
rect 365690 434898 365926 435134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 319610 403718 319846 403954
rect 319610 403398 319846 403634
rect 350330 403718 350566 403954
rect 350330 403398 350566 403634
rect 381050 403718 381286 403954
rect 381050 403398 381286 403634
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 411008 687218 411244 687454
rect 411008 686898 411244 687134
rect 499816 687218 500052 687454
rect 499816 686898 500052 687134
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 410328 655718 410564 655954
rect 410328 655398 410564 655634
rect 500496 655718 500732 655954
rect 500496 655398 500732 655634
rect 411008 651218 411244 651454
rect 411008 650898 411244 651134
rect 499816 651218 500052 651454
rect 499816 650898 500052 651134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 410328 619718 410564 619954
rect 410328 619398 410564 619634
rect 500496 619718 500732 619954
rect 500496 619398 500732 619634
rect 411008 615218 411244 615454
rect 411008 614898 411244 615134
rect 499816 615218 500052 615454
rect 499816 614898 500052 615134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 410328 547718 410564 547954
rect 410328 547398 410564 547634
rect 500496 547718 500732 547954
rect 500496 547398 500732 547634
rect 411008 543218 411244 543454
rect 411008 542898 411244 543134
rect 499816 543218 500052 543454
rect 499816 542898 500052 543134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 410328 511718 410564 511954
rect 410328 511398 410564 511634
rect 500496 511718 500732 511954
rect 500496 511398 500732 511634
rect 411008 507218 411244 507454
rect 411008 506898 411244 507134
rect 499816 507218 500052 507454
rect 499816 506898 500052 507134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 81008 687454
rect 81244 687218 169816 687454
rect 170052 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 191008 687454
rect 191244 687218 279816 687454
rect 280052 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 301008 687454
rect 301244 687218 389816 687454
rect 390052 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 411008 687454
rect 411244 687218 499816 687454
rect 500052 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 81008 687134
rect 81244 686898 169816 687134
rect 170052 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 191008 687134
rect 191244 686898 279816 687134
rect 280052 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 301008 687134
rect 301244 686898 389816 687134
rect 390052 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 411008 687134
rect 411244 686898 499816 687134
rect 500052 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 80328 655954
rect 80564 655718 170496 655954
rect 170732 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 190328 655954
rect 190564 655718 280496 655954
rect 280732 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 300328 655954
rect 300564 655718 390496 655954
rect 390732 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 410328 655954
rect 410564 655718 500496 655954
rect 500732 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 80328 655634
rect 80564 655398 170496 655634
rect 170732 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 190328 655634
rect 190564 655398 280496 655634
rect 280732 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 300328 655634
rect 300564 655398 390496 655634
rect 390732 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 410328 655634
rect 410564 655398 500496 655634
rect 500732 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 81008 651454
rect 81244 651218 169816 651454
rect 170052 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 191008 651454
rect 191244 651218 279816 651454
rect 280052 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 301008 651454
rect 301244 651218 389816 651454
rect 390052 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 411008 651454
rect 411244 651218 499816 651454
rect 500052 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 81008 651134
rect 81244 650898 169816 651134
rect 170052 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 191008 651134
rect 191244 650898 279816 651134
rect 280052 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 301008 651134
rect 301244 650898 389816 651134
rect 390052 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 411008 651134
rect 411244 650898 499816 651134
rect 500052 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 80328 619954
rect 80564 619718 170496 619954
rect 170732 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 190328 619954
rect 190564 619718 280496 619954
rect 280732 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 300328 619954
rect 300564 619718 390496 619954
rect 390732 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 410328 619954
rect 410564 619718 500496 619954
rect 500732 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 80328 619634
rect 80564 619398 170496 619634
rect 170732 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 190328 619634
rect 190564 619398 280496 619634
rect 280732 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 300328 619634
rect 300564 619398 390496 619634
rect 390732 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 410328 619634
rect 410564 619398 500496 619634
rect 500732 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 81008 615454
rect 81244 615218 169816 615454
rect 170052 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 191008 615454
rect 191244 615218 279816 615454
rect 280052 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 301008 615454
rect 301244 615218 389816 615454
rect 390052 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 411008 615454
rect 411244 615218 499816 615454
rect 500052 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 81008 615134
rect 81244 614898 169816 615134
rect 170052 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 191008 615134
rect 191244 614898 279816 615134
rect 280052 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 301008 615134
rect 301244 614898 389816 615134
rect 390052 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 411008 615134
rect 411244 614898 499816 615134
rect 500052 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 80328 547954
rect 80564 547718 170496 547954
rect 170732 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 190328 547954
rect 190564 547718 280496 547954
rect 280732 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 300328 547954
rect 300564 547718 390496 547954
rect 390732 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 410328 547954
rect 410564 547718 500496 547954
rect 500732 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 80328 547634
rect 80564 547398 170496 547634
rect 170732 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 190328 547634
rect 190564 547398 280496 547634
rect 280732 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 300328 547634
rect 300564 547398 390496 547634
rect 390732 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 410328 547634
rect 410564 547398 500496 547634
rect 500732 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 81008 543454
rect 81244 543218 169816 543454
rect 170052 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 191008 543454
rect 191244 543218 279816 543454
rect 280052 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 301008 543454
rect 301244 543218 389816 543454
rect 390052 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 411008 543454
rect 411244 543218 499816 543454
rect 500052 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 81008 543134
rect 81244 542898 169816 543134
rect 170052 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 191008 543134
rect 191244 542898 279816 543134
rect 280052 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 301008 543134
rect 301244 542898 389816 543134
rect 390052 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 411008 543134
rect 411244 542898 499816 543134
rect 500052 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 80328 511954
rect 80564 511718 170496 511954
rect 170732 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 190328 511954
rect 190564 511718 280496 511954
rect 280732 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 300328 511954
rect 300564 511718 390496 511954
rect 390732 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 410328 511954
rect 410564 511718 500496 511954
rect 500732 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 80328 511634
rect 80564 511398 170496 511634
rect 170732 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 190328 511634
rect 190564 511398 280496 511634
rect 280732 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 300328 511634
rect 300564 511398 390496 511634
rect 390732 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 410328 511634
rect 410564 511398 500496 511634
rect 500732 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 81008 507454
rect 81244 507218 169816 507454
rect 170052 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 191008 507454
rect 191244 507218 279816 507454
rect 280052 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 301008 507454
rect 301244 507218 389816 507454
rect 390052 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 411008 507454
rect 411244 507218 499816 507454
rect 500052 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 81008 507134
rect 81244 506898 169816 507134
rect 170052 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 191008 507134
rect 191244 506898 279816 507134
rect 280052 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 301008 507134
rect 301244 506898 389816 507134
rect 390052 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 411008 507134
rect 411244 506898 499816 507134
rect 500052 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 219610 439954
rect 219846 439718 250330 439954
rect 250566 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 319610 439954
rect 319846 439718 350330 439954
rect 350566 439718 381050 439954
rect 381286 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 219610 439634
rect 219846 439398 250330 439634
rect 250566 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 319610 439634
rect 319846 439398 350330 439634
rect 350566 439398 381050 439634
rect 381286 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 304250 435454
rect 304486 435218 334970 435454
rect 335206 435218 365690 435454
rect 365926 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 304250 435134
rect 304486 434898 334970 435134
rect 335206 434898 365690 435134
rect 365926 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 219610 403954
rect 219846 403718 250330 403954
rect 250566 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 319610 403954
rect 319846 403718 350330 403954
rect 350566 403718 381050 403954
rect 381286 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 219610 403634
rect 219846 403398 250330 403634
rect 250566 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 319610 403634
rect 319846 403398 350330 403634
rect 350566 403398 381050 403634
rect 381286 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use cpu  cpu0
timestamp 0
transform 1 0 300000 0 1 400000
box 0 0 84000 56000
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword0
timestamp 0
transform 1 0 80000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword1
timestamp 0
transform 1 0 190000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword2
timestamp 0
transform 1 0 300000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword3
timestamp 0
transform 1 0 410000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword0
timestamp 0
transform 1 0 80000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword1
timestamp 0
transform 1 0 190000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword2
timestamp 0
transform 1 0 300000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword3
timestamp 0
transform 1 0 410000 0 1 490000
box 0 0 91060 89292
use soc_config  mprj
timestamp 0
transform 1 0 200000 0 1 400000
box 1066 0 64898 44000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 691292 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 691292 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 691292 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 691292 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 691292 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 691292 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 691292 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 691292 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 691292 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 691292 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 691292 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 691292 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 691292 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 691292 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 691292 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 691292 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 691292 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 691292 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 691292 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 691292 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 691292 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 691292 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 691292 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 691292 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 446000 231914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 691292 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 446000 267914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 691292 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 691292 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 691292 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 691292 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 691292 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 691292 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 691292 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
