magic
tech sky130B
magscale 1 2
timestamp 1658777287
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 177390 700516 177396 700528
rect 154172 700488 177396 700516
rect 154172 700476 154178 700488
rect 177390 700476 177396 700488
rect 177448 700476 177454 700528
rect 402238 700476 402244 700528
rect 402296 700516 402302 700528
rect 429838 700516 429844 700528
rect 402296 700488 429844 700516
rect 402296 700476 402302 700488
rect 429838 700476 429844 700488
rect 429896 700476 429902 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 173250 700448 173256 700460
rect 137888 700420 173256 700448
rect 137888 700408 137894 700420
rect 173250 700408 173256 700420
rect 173308 700408 173314 700460
rect 188982 700408 188988 700460
rect 189040 700448 189046 700460
rect 202782 700448 202788 700460
rect 189040 700420 202788 700448
rect 189040 700408 189046 700420
rect 202782 700408 202788 700420
rect 202840 700408 202846 700460
rect 298830 700408 298836 700460
rect 298888 700448 298894 700460
rect 332502 700448 332508 700460
rect 298888 700420 332508 700448
rect 298888 700408 298894 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 402330 700408 402336 700460
rect 402388 700448 402394 700460
rect 462314 700448 462320 700460
rect 402388 700420 462320 700448
rect 402388 700408 402394 700420
rect 462314 700408 462320 700420
rect 462372 700408 462378 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 33778 700380 33784 700392
rect 24360 700352 33784 700380
rect 24360 700340 24366 700352
rect 33778 700340 33784 700352
rect 33836 700340 33842 700392
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 51718 700380 51724 700392
rect 40552 700352 51724 700380
rect 40552 700340 40558 700352
rect 51718 700340 51724 700352
rect 51776 700340 51782 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 177298 700380 177304 700392
rect 105504 700352 177304 700380
rect 105504 700340 105510 700352
rect 177298 700340 177304 700352
rect 177356 700340 177362 700392
rect 189994 700340 190000 700392
rect 190052 700380 190058 700392
rect 218974 700380 218980 700392
rect 190052 700352 218980 700380
rect 190052 700340 190058 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 290550 700340 290556 700392
rect 290608 700380 290614 700392
rect 348786 700380 348792 700392
rect 290608 700352 348792 700380
rect 290608 700340 290614 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 392578 700340 392584 700392
rect 392636 700380 392642 700392
rect 478506 700380 478512 700392
rect 392636 700352 478512 700380
rect 392636 700340 392642 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 55858 700312 55864 700324
rect 8168 700284 55864 700312
rect 8168 700272 8174 700284
rect 55858 700272 55864 700284
rect 55916 700272 55922 700324
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 171778 700312 171784 700324
rect 89220 700284 171784 700312
rect 89220 700272 89226 700284
rect 171778 700272 171784 700284
rect 171836 700272 171842 700324
rect 189902 700272 189908 700324
rect 189960 700312 189966 700324
rect 235166 700312 235172 700324
rect 189960 700284 235172 700312
rect 189960 700272 189966 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 281534 700312 281540 700324
rect 267700 700284 281540 700312
rect 267700 700272 267706 700284
rect 281534 700272 281540 700284
rect 281592 700272 281598 700324
rect 294598 700272 294604 700324
rect 294656 700312 294662 700324
rect 364978 700312 364984 700324
rect 294656 700284 364984 700312
rect 294656 700272 294662 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 393958 700272 393964 700324
rect 394016 700312 394022 700324
rect 494790 700312 494796 700324
rect 394016 700284 494796 700312
rect 394016 700272 394022 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 505738 700272 505744 700324
rect 505796 700312 505802 700324
rect 559650 700312 559656 700324
rect 505796 700284 559656 700312
rect 505796 700272 505802 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 173158 699700 173164 699712
rect 170364 699672 173164 699700
rect 170364 699660 170370 699672
rect 173158 699660 173164 699672
rect 173216 699660 173222 699712
rect 298738 699660 298744 699712
rect 298796 699700 298802 699712
rect 300118 699700 300124 699712
rect 298796 699672 300124 699700
rect 298796 699660 298802 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 409138 699660 409144 699712
rect 409196 699700 409202 699712
rect 413646 699700 413652 699712
rect 409196 699672 413652 699700
rect 409196 699660 409202 699672
rect 413646 699660 413652 699672
rect 413704 699660 413710 699712
rect 290458 696940 290464 696992
rect 290516 696980 290522 696992
rect 580166 696980 580172 696992
rect 290516 696952 580172 696980
rect 290516 696940 290522 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 15838 683176 15844 683188
rect 3476 683148 15844 683176
rect 3476 683136 3482 683148
rect 15838 683136 15844 683148
rect 15896 683136 15902 683188
rect 533338 683136 533344 683188
rect 533396 683176 533402 683188
rect 580166 683176 580172 683188
rect 533396 683148 580172 683176
rect 533396 683136 533402 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 37918 670732 37924 670744
rect 3568 670704 37924 670732
rect 3568 670692 3574 670704
rect 37918 670692 37924 670704
rect 37976 670692 37982 670744
rect 502978 670692 502984 670744
rect 503036 670732 503042 670744
rect 580166 670732 580172 670744
rect 503036 670704 580172 670732
rect 503036 670692 503042 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4798 656996 4804 657008
rect 2832 656968 4804 656996
rect 2832 656956 2838 656968
rect 4798 656956 4804 656968
rect 4856 656956 4862 657008
rect 503070 643084 503076 643136
rect 503128 643124 503134 643136
rect 580166 643124 580172 643136
rect 503128 643096 580172 643124
rect 503128 643084 503134 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 51810 632108 51816 632120
rect 3476 632080 51816 632108
rect 3476 632068 3482 632080
rect 51810 632068 51816 632080
rect 51868 632068 51874 632120
rect 523678 630640 523684 630692
rect 523736 630680 523742 630692
rect 580166 630680 580172 630692
rect 523736 630652 580172 630680
rect 523736 630640 523742 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 503162 616836 503168 616888
rect 503220 616876 503226 616888
rect 580166 616876 580172 616888
rect 503220 616848 580172 616876
rect 503220 616836 503226 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3142 605888 3148 605940
rect 3200 605928 3206 605940
rect 6178 605928 6184 605940
rect 3200 605900 6184 605928
rect 3200 605888 3206 605900
rect 6178 605888 6184 605900
rect 6236 605888 6242 605940
rect 407758 600244 407764 600296
rect 407816 600284 407822 600296
rect 407942 600284 407948 600296
rect 407816 600256 407948 600284
rect 407816 600244 407822 600256
rect 407942 600244 407948 600256
rect 408000 600244 408006 600296
rect 78122 599972 78128 600024
rect 78180 600012 78186 600024
rect 187234 600012 187240 600024
rect 78180 599984 187240 600012
rect 78180 599972 78186 599984
rect 187234 599972 187240 599984
rect 187292 599972 187298 600024
rect 297818 599972 297824 600024
rect 297876 600012 297882 600024
rect 408218 600012 408224 600024
rect 297876 599984 408224 600012
rect 297876 599972 297882 599984
rect 408218 599972 408224 599984
rect 408276 599972 408282 600024
rect 78030 599904 78036 599956
rect 78088 599944 78094 599956
rect 187142 599944 187148 599956
rect 78088 599916 187148 599944
rect 78088 599904 78094 599916
rect 187142 599904 187148 599916
rect 187200 599904 187206 599956
rect 78214 599836 78220 599888
rect 78272 599876 78278 599888
rect 187326 599876 187332 599888
rect 78272 599848 187332 599876
rect 78272 599836 78278 599848
rect 187326 599836 187332 599848
rect 187384 599836 187390 599888
rect 78582 599768 78588 599820
rect 78640 599808 78646 599820
rect 186590 599808 186596 599820
rect 78640 599780 186596 599808
rect 78640 599768 78646 599780
rect 186590 599768 186596 599780
rect 186648 599768 186654 599820
rect 297358 599768 297364 599820
rect 297416 599808 297422 599820
rect 297818 599808 297824 599820
rect 297416 599780 297824 599808
rect 297416 599768 297422 599780
rect 297818 599768 297824 599780
rect 297876 599768 297882 599820
rect 78398 599700 78404 599752
rect 78456 599740 78462 599752
rect 187050 599740 187056 599752
rect 78456 599712 187056 599740
rect 78456 599700 78462 599712
rect 187050 599700 187056 599712
rect 187108 599700 187114 599752
rect 78490 599632 78496 599684
rect 78548 599672 78554 599684
rect 186866 599672 186872 599684
rect 78548 599644 186872 599672
rect 78548 599632 78554 599644
rect 186866 599632 186872 599644
rect 186924 599632 186930 599684
rect 297910 599564 297916 599616
rect 297968 599604 297974 599616
rect 407758 599604 407764 599616
rect 297968 599576 407764 599604
rect 297968 599564 297974 599576
rect 407758 599564 407764 599576
rect 407816 599564 407822 599616
rect 297266 599360 297272 599412
rect 297324 599400 297330 599412
rect 297910 599400 297916 599412
rect 297324 599372 297916 599400
rect 297324 599360 297330 599372
rect 297910 599360 297916 599372
rect 297968 599360 297974 599412
rect 297450 598884 297456 598936
rect 297508 598924 297514 598936
rect 407574 598924 407580 598936
rect 297508 598896 407580 598924
rect 297508 598884 297514 598896
rect 407574 598884 407580 598896
rect 407632 598884 407638 598936
rect 297542 598816 297548 598868
rect 297600 598856 297606 598868
rect 407390 598856 407396 598868
rect 297600 598828 407396 598856
rect 297600 598816 297606 598828
rect 407390 598816 407396 598828
rect 407448 598816 407454 598868
rect 297174 598272 297180 598324
rect 297232 598312 297238 598324
rect 298002 598312 298008 598324
rect 297232 598284 298008 598312
rect 297232 598272 297238 598284
rect 298002 598272 298008 598284
rect 298060 598312 298066 598324
rect 298060 598284 306374 598312
rect 298060 598272 298066 598284
rect 306346 598244 306374 598284
rect 407482 598244 407488 598256
rect 306346 598216 407488 598244
rect 407482 598204 407488 598216
rect 407540 598204 407546 598256
rect 115842 597524 115848 597576
rect 115900 597564 115906 597576
rect 225506 597564 225512 597576
rect 115900 597536 225512 597564
rect 115900 597524 115906 597536
rect 225506 597524 225512 597536
rect 225564 597564 225570 597576
rect 282362 597564 282368 597576
rect 225564 597536 282368 597564
rect 225564 597524 225570 597536
rect 282362 597524 282368 597536
rect 282420 597564 282426 597576
rect 335354 597564 335360 597576
rect 282420 597536 335360 597564
rect 282420 597524 282426 597536
rect 335354 597524 335360 597536
rect 335412 597564 335418 597576
rect 444374 597564 444380 597576
rect 335412 597536 444380 597564
rect 335412 597524 335418 597536
rect 444374 597524 444380 597536
rect 444432 597524 444438 597576
rect 126882 597456 126888 597508
rect 126940 597496 126946 597508
rect 234614 597496 234620 597508
rect 126940 597468 234620 597496
rect 126940 597456 126946 597468
rect 234614 597456 234620 597468
rect 234672 597456 234678 597508
rect 326154 597456 326160 597508
rect 326212 597496 326218 597508
rect 434714 597496 434720 597508
rect 326212 597468 434720 597496
rect 326212 597456 326218 597468
rect 434714 597456 434720 597468
rect 434772 597456 434778 597508
rect 136542 597388 136548 597440
rect 136600 597428 136606 597440
rect 245470 597428 245476 597440
rect 136600 597400 245476 597428
rect 136600 597388 136606 597400
rect 245470 597388 245476 597400
rect 245528 597428 245534 597440
rect 245528 597400 248414 597428
rect 245528 597388 245534 597400
rect 111702 597320 111708 597372
rect 111760 597360 111766 597372
rect 219434 597360 219440 597372
rect 111760 597332 219440 597360
rect 111760 597320 111766 597332
rect 219434 597320 219440 597332
rect 219492 597360 219498 597372
rect 220722 597360 220728 597372
rect 219492 597332 220728 597360
rect 219492 597320 219498 597332
rect 220722 597320 220728 597332
rect 220780 597320 220786 597372
rect 103146 597252 103152 597304
rect 103204 597292 103210 597304
rect 212350 597292 212356 597304
rect 103204 597264 212356 597292
rect 103204 597252 103210 597264
rect 212350 597252 212356 597264
rect 212408 597252 212414 597304
rect 140682 597184 140688 597236
rect 140740 597224 140746 597236
rect 140740 597196 243584 597224
rect 140740 597184 140746 597196
rect 131022 597116 131028 597168
rect 131080 597156 131086 597168
rect 131080 597128 238754 597156
rect 131080 597116 131086 597128
rect 106182 597048 106188 597100
rect 106240 597088 106246 597100
rect 215294 597088 215300 597100
rect 106240 597060 215300 597088
rect 106240 597048 106246 597060
rect 215294 597048 215300 597060
rect 215352 597048 215358 597100
rect 121362 596980 121368 597032
rect 121420 597020 121426 597032
rect 121420 596992 219434 597020
rect 121420 596980 121426 596992
rect 100662 596912 100668 596964
rect 100720 596952 100726 596964
rect 209958 596952 209964 596964
rect 100720 596924 209964 596952
rect 100720 596912 100726 596924
rect 209958 596912 209964 596924
rect 210016 596952 210022 596964
rect 211062 596952 211068 596964
rect 210016 596924 211068 596952
rect 210016 596912 210022 596924
rect 211062 596912 211068 596924
rect 211120 596912 211126 596964
rect 103422 596844 103428 596896
rect 103480 596884 103486 596896
rect 213822 596884 213828 596896
rect 103480 596856 213828 596884
rect 103480 596844 103486 596856
rect 213822 596844 213828 596856
rect 213880 596844 213886 596896
rect 104802 596776 104808 596828
rect 104860 596816 104866 596828
rect 214834 596816 214840 596828
rect 104860 596788 214840 596816
rect 104860 596776 104866 596788
rect 214834 596776 214840 596788
rect 214892 596776 214898 596828
rect 219406 596816 219434 596992
rect 238726 596952 238754 597128
rect 243556 597088 243584 597196
rect 248386 597156 248414 597400
rect 281626 597388 281632 597440
rect 281684 597428 281690 597440
rect 350442 597428 350448 597440
rect 281684 597400 350448 597428
rect 281684 597388 281690 597400
rect 350442 597388 350448 597400
rect 350500 597428 350506 597440
rect 459554 597428 459560 597440
rect 350500 597400 459560 597428
rect 350500 597388 350506 597400
rect 459554 597388 459560 597400
rect 459612 597388 459618 597440
rect 330386 597320 330392 597372
rect 330444 597360 330450 597372
rect 440234 597360 440240 597372
rect 330444 597332 440240 597360
rect 330444 597320 330450 597332
rect 440234 597320 440240 597332
rect 440292 597320 440298 597372
rect 281718 597252 281724 597304
rect 281776 597292 281782 597304
rect 345658 597292 345664 597304
rect 281776 597264 345664 597292
rect 281776 597252 281782 597264
rect 345658 597252 345664 597264
rect 345716 597292 345722 597304
rect 455414 597292 455420 597304
rect 345716 597264 455420 597292
rect 345716 597252 345722 597264
rect 455414 597252 455420 597264
rect 455472 597252 455478 597304
rect 282178 597184 282184 597236
rect 282236 597224 282242 597236
rect 340506 597224 340512 597236
rect 282236 597196 340512 597224
rect 282236 597184 282242 597196
rect 340506 597184 340512 597196
rect 340564 597224 340570 597236
rect 449894 597224 449900 597236
rect 340564 597196 449900 597224
rect 340564 597184 340570 597196
rect 449894 597184 449900 597196
rect 449952 597184 449958 597236
rect 282086 597156 282092 597168
rect 248386 597128 282092 597156
rect 282086 597116 282092 597128
rect 282144 597116 282150 597168
rect 323394 597156 323400 597168
rect 316006 597128 323400 597156
rect 250530 597088 250536 597100
rect 243556 597060 250536 597088
rect 250530 597048 250536 597060
rect 250588 597088 250594 597100
rect 250588 597060 277394 597088
rect 250588 597048 250594 597060
rect 277366 597020 277394 597060
rect 284294 597048 284300 597100
rect 284352 597088 284358 597100
rect 316006 597088 316034 597128
rect 323394 597116 323400 597128
rect 323452 597156 323458 597168
rect 433334 597156 433340 597168
rect 323452 597128 433340 597156
rect 323452 597116 323458 597128
rect 433334 597116 433340 597128
rect 433392 597116 433398 597168
rect 284352 597060 316034 597088
rect 284352 597048 284358 597060
rect 324314 597048 324320 597100
rect 324372 597088 324378 597100
rect 324774 597088 324780 597100
rect 324372 597060 324780 597088
rect 324372 597048 324378 597060
rect 324774 597048 324780 597060
rect 324832 597088 324838 597100
rect 434714 597088 434720 597100
rect 324832 597060 434720 597088
rect 324832 597048 324838 597060
rect 434714 597048 434720 597060
rect 434772 597048 434778 597100
rect 281902 597020 281908 597032
rect 277366 596992 281908 597020
rect 281902 596980 281908 596992
rect 281960 597020 281966 597032
rect 360562 597020 360568 597032
rect 281960 596992 360568 597020
rect 281960 596980 281966 596992
rect 360562 596980 360568 596992
rect 360620 597020 360626 597032
rect 360620 596992 364334 597020
rect 360620 596980 360626 596992
rect 240502 596952 240508 596964
rect 238726 596924 240508 596952
rect 240502 596912 240508 596924
rect 240560 596952 240566 596964
rect 281626 596952 281632 596964
rect 240560 596924 281632 596952
rect 240560 596912 240566 596924
rect 281626 596912 281632 596924
rect 281684 596912 281690 596964
rect 281994 596912 282000 596964
rect 282052 596952 282058 596964
rect 284662 596952 284668 596964
rect 282052 596924 284668 596952
rect 282052 596912 282058 596924
rect 284662 596912 284668 596924
rect 284720 596912 284726 596964
rect 299382 596912 299388 596964
rect 299440 596952 299446 596964
rect 314654 596952 314660 596964
rect 299440 596924 314660 596952
rect 299440 596912 299446 596924
rect 314654 596912 314660 596924
rect 314712 596912 314718 596964
rect 364306 596952 364334 596992
rect 470594 596952 470600 596964
rect 364306 596924 470600 596952
rect 470594 596912 470600 596924
rect 470652 596912 470658 596964
rect 234614 596844 234620 596896
rect 234672 596884 234678 596896
rect 281718 596884 281724 596896
rect 234672 596856 281724 596884
rect 234672 596844 234678 596856
rect 281718 596844 281724 596856
rect 281776 596844 281782 596896
rect 282270 596844 282276 596896
rect 282328 596884 282334 596896
rect 319990 596884 319996 596896
rect 282328 596856 319996 596884
rect 282328 596844 282334 596856
rect 319990 596844 319996 596856
rect 320048 596884 320054 596896
rect 429194 596884 429200 596896
rect 320048 596856 429200 596884
rect 320048 596844 320054 596856
rect 429194 596844 429200 596856
rect 429252 596844 429258 596896
rect 230658 596816 230664 596828
rect 219406 596788 230664 596816
rect 230658 596776 230664 596788
rect 230716 596816 230722 596828
rect 282178 596816 282184 596828
rect 230716 596788 282184 596816
rect 230716 596776 230722 596788
rect 282178 596776 282184 596788
rect 282236 596776 282242 596828
rect 284938 596776 284944 596828
rect 284996 596816 285002 596828
rect 322290 596816 322296 596828
rect 284996 596788 322296 596816
rect 284996 596776 285002 596788
rect 322290 596776 322296 596788
rect 322348 596816 322354 596828
rect 431954 596816 431960 596828
rect 322348 596788 431960 596816
rect 322348 596776 322354 596788
rect 431954 596776 431960 596788
rect 432012 596776 432018 596828
rect 220722 596708 220728 596760
rect 220780 596748 220786 596760
rect 280982 596748 280988 596760
rect 220780 596720 280988 596748
rect 220780 596708 220786 596720
rect 280982 596708 280988 596720
rect 281040 596748 281046 596760
rect 330386 596748 330392 596760
rect 281040 596720 330392 596748
rect 281040 596708 281046 596720
rect 330386 596708 330392 596720
rect 330444 596708 330450 596760
rect 354674 596748 354680 596760
rect 354646 596708 354680 596748
rect 354732 596748 354738 596760
rect 465074 596748 465080 596760
rect 354732 596720 465080 596748
rect 354732 596708 354738 596720
rect 465074 596708 465080 596720
rect 465132 596708 465138 596760
rect 215294 596640 215300 596692
rect 215352 596680 215358 596692
rect 284570 596680 284576 596692
rect 215352 596652 284576 596680
rect 215352 596640 215358 596652
rect 284570 596640 284576 596652
rect 284628 596640 284634 596692
rect 214834 596572 214840 596624
rect 214892 596612 214898 596624
rect 284478 596612 284484 596624
rect 214892 596584 284484 596612
rect 214892 596572 214898 596584
rect 284478 596572 284484 596584
rect 284536 596612 284542 596624
rect 324314 596612 324320 596624
rect 284536 596584 324320 596612
rect 284536 596572 284542 596584
rect 324314 596572 324320 596584
rect 324372 596572 324378 596624
rect 213822 596504 213828 596556
rect 213880 596544 213886 596556
rect 284294 596544 284300 596556
rect 213880 596516 284300 596544
rect 213880 596504 213886 596516
rect 284294 596504 284300 596516
rect 284352 596504 284358 596556
rect 284570 596504 284576 596556
rect 284628 596544 284634 596556
rect 326154 596544 326160 596556
rect 284628 596516 326160 596544
rect 284628 596504 284634 596516
rect 326154 596504 326160 596516
rect 326212 596504 326218 596556
rect 212442 596436 212448 596488
rect 212500 596476 212506 596488
rect 284386 596476 284392 596488
rect 212500 596448 284392 596476
rect 212500 596436 212506 596448
rect 284386 596436 284392 596448
rect 284444 596436 284450 596488
rect 211062 596368 211068 596420
rect 211120 596408 211126 596420
rect 282270 596408 282276 596420
rect 211120 596380 282276 596408
rect 211120 596368 211126 596380
rect 282270 596368 282276 596380
rect 282328 596368 282334 596420
rect 354646 596408 354674 596708
rect 287026 596380 354674 596408
rect 79778 596300 79784 596352
rect 79836 596340 79842 596352
rect 92474 596340 92480 596352
rect 79836 596312 92480 596340
rect 79836 596300 79842 596312
rect 92474 596300 92480 596312
rect 92532 596300 92538 596352
rect 188706 596300 188712 596352
rect 188764 596340 188770 596352
rect 202874 596340 202880 596352
rect 188764 596312 202880 596340
rect 188764 596300 188770 596312
rect 202874 596300 202880 596312
rect 202932 596300 202938 596352
rect 209038 596300 209044 596352
rect 209096 596340 209102 596352
rect 281994 596340 282000 596352
rect 209096 596312 282000 596340
rect 209096 596300 209102 596312
rect 281994 596300 282000 596312
rect 282052 596300 282058 596352
rect 282086 596300 282092 596352
rect 282144 596340 282150 596352
rect 287026 596340 287054 596380
rect 282144 596312 287054 596340
rect 282144 596300 282150 596312
rect 408218 596300 408224 596352
rect 408276 596340 408282 596352
rect 422570 596340 422576 596352
rect 408276 596312 422576 596340
rect 408276 596300 408282 596312
rect 422570 596300 422576 596312
rect 422628 596300 422634 596352
rect 79870 596232 79876 596284
rect 79928 596272 79934 596284
rect 94038 596272 94044 596284
rect 79928 596244 94044 596272
rect 79928 596232 79934 596244
rect 94038 596232 94044 596244
rect 94096 596232 94102 596284
rect 188890 596232 188896 596284
rect 188948 596272 188954 596284
rect 204346 596272 204352 596284
rect 188948 596244 204352 596272
rect 188948 596232 188954 596244
rect 204346 596232 204352 596244
rect 204404 596232 204410 596284
rect 207658 596232 207664 596284
rect 207716 596272 207722 596284
rect 284754 596272 284760 596284
rect 207716 596244 284760 596272
rect 207716 596232 207722 596244
rect 284754 596232 284760 596244
rect 284812 596232 284818 596284
rect 299290 596232 299296 596284
rect 299348 596272 299354 596284
rect 311894 596272 311900 596284
rect 299348 596244 311900 596272
rect 299348 596232 299354 596244
rect 311894 596232 311900 596244
rect 311952 596232 311958 596284
rect 407942 596232 407948 596284
rect 408000 596272 408006 596284
rect 423674 596272 423680 596284
rect 408000 596244 423680 596272
rect 408000 596232 408006 596244
rect 423674 596232 423680 596244
rect 423732 596232 423738 596284
rect 79962 596164 79968 596216
rect 80020 596204 80026 596216
rect 95234 596204 95240 596216
rect 80020 596176 95240 596204
rect 80020 596164 80026 596176
rect 95234 596164 95240 596176
rect 95292 596164 95298 596216
rect 188798 596164 188804 596216
rect 188856 596204 188862 596216
rect 204254 596204 204260 596216
rect 188856 596176 204260 596204
rect 188856 596164 188862 596176
rect 204254 596164 204260 596176
rect 204312 596164 204318 596216
rect 212350 596164 212356 596216
rect 212408 596204 212414 596216
rect 284938 596204 284944 596216
rect 212408 596176 284944 596204
rect 212408 596164 212414 596176
rect 284938 596164 284944 596176
rect 284996 596164 285002 596216
rect 299198 596164 299204 596216
rect 299256 596204 299262 596216
rect 313274 596204 313280 596216
rect 299256 596176 313280 596204
rect 299256 596164 299262 596176
rect 313274 596164 313280 596176
rect 313332 596164 313338 596216
rect 407758 596164 407764 596216
rect 407816 596204 407822 596216
rect 425054 596204 425060 596216
rect 407816 596176 425060 596204
rect 407816 596164 407822 596176
rect 425054 596164 425060 596176
rect 425112 596164 425118 596216
rect 281626 591336 281632 591388
rect 281684 591376 281690 591388
rect 281994 591376 282000 591388
rect 281684 591348 282000 591376
rect 281684 591336 281690 591348
rect 281994 591336 282000 591348
rect 282052 591336 282058 591388
rect 281626 591200 281632 591252
rect 281684 591240 281690 591252
rect 282362 591240 282368 591252
rect 281684 591212 282368 591240
rect 281684 591200 281690 591212
rect 282362 591200 282368 591212
rect 282420 591200 282426 591252
rect 283558 590656 283564 590708
rect 283616 590696 283622 590708
rect 579798 590696 579804 590708
rect 283616 590668 579804 590696
rect 283616 590656 283622 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 78306 584400 78312 584452
rect 78364 584440 78370 584452
rect 186682 584440 186688 584452
rect 78364 584412 186688 584440
rect 78364 584400 78370 584412
rect 186682 584400 186688 584412
rect 186740 584400 186746 584452
rect 2774 579912 2780 579964
rect 2832 579952 2838 579964
rect 4890 579952 4896 579964
rect 2832 579924 4896 579952
rect 2832 579912 2838 579924
rect 4890 579912 4896 579924
rect 4948 579912 4954 579964
rect 501598 563048 501604 563100
rect 501656 563088 501662 563100
rect 580166 563088 580172 563100
rect 501656 563060 580172 563088
rect 501656 563048 501662 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553528 3332 553580
rect 3384 553568 3390 553580
rect 7558 553568 7564 553580
rect 3384 553540 7564 553568
rect 3384 553528 3390 553540
rect 7558 553528 7564 553540
rect 7616 553528 7622 553580
rect 515398 536800 515404 536852
rect 515456 536840 515462 536852
rect 579890 536840 579896 536852
rect 515456 536812 579896 536840
rect 515456 536800 515462 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2774 527212 2780 527264
rect 2832 527252 2838 527264
rect 4982 527252 4988 527264
rect 2832 527224 4988 527252
rect 2832 527212 2838 527224
rect 4982 527212 4988 527224
rect 5040 527212 5046 527264
rect 284938 526396 284944 526448
rect 284996 526436 285002 526448
rect 297174 526436 297180 526448
rect 284996 526408 297180 526436
rect 284996 526396 285002 526408
rect 297174 526396 297180 526408
rect 297232 526436 297238 526448
rect 297726 526436 297732 526448
rect 297232 526408 297732 526436
rect 297232 526396 297238 526408
rect 297726 526396 297732 526408
rect 297784 526396 297790 526448
rect 294690 525920 294696 525972
rect 294748 525960 294754 525972
rect 297266 525960 297272 525972
rect 294748 525932 297272 525960
rect 294748 525920 294754 525932
rect 297266 525920 297272 525932
rect 297324 525960 297330 525972
rect 298002 525960 298008 525972
rect 297324 525932 298008 525960
rect 297324 525920 297330 525932
rect 298002 525920 298008 525932
rect 298060 525920 298066 525972
rect 186866 525852 186872 525904
rect 186924 525892 186930 525904
rect 187694 525892 187700 525904
rect 186924 525864 187700 525892
rect 186924 525852 186930 525864
rect 187694 525852 187700 525864
rect 187752 525852 187758 525904
rect 519538 524424 519544 524476
rect 519596 524464 519602 524476
rect 580166 524464 580172 524476
rect 519596 524436 580172 524464
rect 519596 524424 519602 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 285582 523744 285588 523796
rect 285640 523784 285646 523796
rect 297358 523784 297364 523796
rect 285640 523756 297364 523784
rect 285640 523744 285646 523756
rect 297358 523744 297364 523756
rect 297416 523784 297422 523796
rect 298002 523784 298008 523796
rect 297416 523756 298008 523784
rect 297416 523744 297422 523756
rect 298002 523744 298008 523756
rect 298060 523744 298066 523796
rect 284202 523676 284208 523728
rect 284260 523716 284266 523728
rect 297634 523716 297640 523728
rect 284260 523688 297640 523716
rect 284260 523676 284266 523688
rect 297634 523676 297640 523688
rect 297692 523716 297698 523728
rect 297910 523716 297916 523728
rect 297692 523688 297916 523716
rect 297692 523676 297698 523688
rect 297910 523676 297916 523688
rect 297968 523676 297974 523728
rect 187510 521568 187516 521620
rect 187568 521608 187574 521620
rect 188154 521608 188160 521620
rect 187568 521580 188160 521608
rect 187568 521568 187574 521580
rect 188154 521568 188160 521580
rect 188212 521568 188218 521620
rect 284110 520956 284116 521008
rect 284168 520996 284174 521008
rect 297450 520996 297456 521008
rect 284168 520968 297456 520996
rect 284168 520956 284174 520968
rect 297450 520956 297456 520968
rect 297508 520956 297514 521008
rect 284018 520888 284024 520940
rect 284076 520928 284082 520940
rect 297818 520928 297824 520940
rect 284076 520900 297824 520928
rect 284076 520888 284082 520900
rect 297818 520888 297824 520900
rect 297876 520888 297882 520940
rect 187142 518372 187148 518424
rect 187200 518412 187206 518424
rect 188062 518412 188068 518424
rect 187200 518384 188068 518412
rect 187200 518372 187206 518384
rect 188062 518372 188068 518384
rect 188120 518372 188126 518424
rect 282822 518168 282828 518220
rect 282880 518208 282886 518220
rect 297542 518208 297548 518220
rect 282880 518180 297548 518208
rect 282880 518168 282886 518180
rect 297542 518168 297548 518180
rect 297600 518168 297606 518220
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 14458 514808 14464 514820
rect 3384 514780 14464 514808
rect 3384 514768 3390 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 549898 510620 549904 510672
rect 549956 510660 549962 510672
rect 580166 510660 580172 510672
rect 549956 510632 580172 510660
rect 549956 510620 549962 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 15930 501004 15936 501016
rect 3384 500976 15936 501004
rect 3384 500964 3390 500976
rect 15930 500964 15936 500976
rect 15988 500964 15994 501016
rect 78122 489812 78128 489864
rect 78180 489852 78186 489864
rect 187970 489852 187976 489864
rect 78180 489824 187976 489852
rect 78180 489812 78186 489824
rect 187970 489812 187976 489824
rect 188028 489812 188034 489864
rect 408126 489852 408132 489864
rect 284036 489824 408132 489852
rect 284036 489796 284064 489824
rect 408126 489812 408132 489824
rect 408184 489812 408190 489864
rect 78030 489744 78036 489796
rect 78088 489784 78094 489796
rect 188062 489784 188068 489796
rect 78088 489756 188068 489784
rect 78088 489744 78094 489756
rect 188062 489744 188068 489756
rect 188120 489744 188126 489796
rect 284018 489744 284024 489796
rect 284076 489744 284082 489796
rect 284202 489744 284208 489796
rect 284260 489784 284266 489796
rect 407666 489784 407672 489796
rect 284260 489756 407672 489784
rect 284260 489744 284266 489756
rect 407666 489744 407672 489756
rect 407724 489744 407730 489796
rect 77754 489676 77760 489728
rect 77812 489716 77818 489728
rect 188154 489716 188160 489728
rect 77812 489688 188160 489716
rect 77812 489676 77818 489688
rect 188154 489676 188160 489688
rect 188212 489676 188218 489728
rect 284110 489676 284116 489728
rect 284168 489716 284174 489728
rect 407574 489716 407580 489728
rect 284168 489688 407580 489716
rect 284168 489676 284174 489688
rect 407574 489676 407580 489688
rect 407632 489676 407638 489728
rect 78306 489608 78312 489660
rect 78364 489648 78370 489660
rect 188338 489648 188344 489660
rect 78364 489620 188344 489648
rect 78364 489608 78370 489620
rect 188338 489608 188344 489620
rect 188396 489608 188402 489660
rect 297910 489608 297916 489660
rect 297968 489648 297974 489660
rect 408402 489648 408408 489660
rect 297968 489620 408408 489648
rect 297968 489608 297974 489620
rect 408402 489608 408408 489620
rect 408460 489608 408466 489660
rect 77570 489540 77576 489592
rect 77628 489580 77634 489592
rect 187786 489580 187792 489592
rect 77628 489552 187792 489580
rect 77628 489540 77634 489552
rect 187786 489540 187792 489552
rect 187844 489540 187850 489592
rect 297818 489540 297824 489592
rect 297876 489580 297882 489592
rect 407850 489580 407856 489592
rect 297876 489552 407856 489580
rect 297876 489540 297882 489552
rect 407850 489540 407856 489552
rect 407908 489540 407914 489592
rect 78490 489472 78496 489524
rect 78548 489512 78554 489524
rect 187694 489512 187700 489524
rect 78548 489484 187700 489512
rect 78548 489472 78554 489484
rect 187694 489472 187700 489484
rect 187752 489472 187758 489524
rect 77662 489404 77668 489456
rect 77720 489444 77726 489456
rect 187050 489444 187056 489456
rect 77720 489416 187056 489444
rect 77720 489404 77726 489416
rect 187050 489404 187056 489416
rect 187108 489404 187114 489456
rect 78582 489336 78588 489388
rect 78640 489376 78646 489388
rect 186958 489376 186964 489388
rect 78640 489348 186964 489376
rect 78640 489336 78646 489348
rect 186958 489336 186964 489348
rect 187016 489336 187022 489388
rect 188338 489132 188344 489184
rect 188396 489172 188402 489184
rect 240778 489172 240784 489184
rect 188396 489144 240784 489172
rect 188396 489132 188402 489144
rect 240778 489132 240784 489144
rect 240836 489132 240842 489184
rect 187970 488860 187976 488912
rect 188028 488900 188034 488912
rect 188614 488900 188620 488912
rect 188028 488872 188620 488900
rect 188028 488860 188034 488872
rect 188614 488860 188620 488872
rect 188672 488860 188678 488912
rect 110506 488792 110512 488844
rect 110564 488832 110570 488844
rect 220722 488832 220728 488844
rect 110564 488804 220728 488832
rect 110564 488792 110570 488804
rect 220722 488792 220728 488804
rect 220780 488792 220786 488844
rect 187786 488724 187792 488776
rect 187844 488764 187850 488776
rect 188246 488764 188252 488776
rect 187844 488736 188252 488764
rect 187844 488724 187850 488736
rect 188246 488724 188252 488736
rect 188304 488724 188310 488776
rect 215294 488724 215300 488776
rect 215352 488764 215358 488776
rect 242894 488764 242900 488776
rect 215352 488736 242900 488764
rect 215352 488724 215358 488736
rect 242894 488724 242900 488736
rect 242952 488764 242958 488776
rect 325326 488764 325332 488776
rect 242952 488736 325332 488764
rect 242952 488724 242958 488736
rect 325326 488724 325332 488736
rect 325384 488764 325390 488776
rect 325384 488736 325694 488764
rect 325384 488724 325390 488736
rect 120626 488656 120632 488708
rect 120684 488696 120690 488708
rect 230474 488696 230480 488708
rect 120684 488668 230480 488696
rect 120684 488656 120690 488668
rect 230474 488656 230480 488668
rect 230532 488696 230538 488708
rect 231762 488696 231768 488708
rect 230532 488668 231768 488696
rect 230532 488656 230538 488668
rect 231762 488656 231768 488668
rect 231820 488656 231826 488708
rect 283650 488656 283656 488708
rect 283708 488696 283714 488708
rect 284202 488696 284208 488708
rect 283708 488668 284208 488696
rect 283708 488656 283714 488668
rect 284202 488656 284208 488668
rect 284260 488656 284266 488708
rect 297358 488656 297364 488708
rect 297416 488696 297422 488708
rect 297818 488696 297824 488708
rect 297416 488668 297824 488696
rect 297416 488656 297422 488668
rect 297818 488656 297824 488668
rect 297876 488656 297882 488708
rect 325666 488696 325694 488736
rect 336642 488724 336648 488776
rect 336700 488764 336706 488776
rect 444374 488764 444380 488776
rect 336700 488736 444380 488764
rect 336700 488724 336706 488736
rect 444374 488724 444380 488736
rect 444432 488724 444438 488776
rect 434714 488696 434720 488708
rect 325666 488668 434720 488696
rect 434714 488656 434720 488668
rect 434772 488656 434778 488708
rect 115658 488588 115664 488640
rect 115716 488628 115722 488640
rect 226242 488628 226248 488640
rect 115716 488600 226248 488628
rect 115716 488588 115722 488600
rect 226242 488588 226248 488600
rect 226300 488628 226306 488640
rect 335446 488628 335452 488640
rect 226300 488600 335452 488628
rect 226300 488588 226306 488600
rect 335446 488588 335452 488600
rect 335504 488628 335510 488640
rect 336642 488628 336648 488640
rect 335504 488600 336648 488628
rect 335504 488588 335510 488600
rect 336642 488588 336648 488600
rect 336700 488588 336706 488640
rect 340598 488588 340604 488640
rect 340656 488628 340662 488640
rect 449894 488628 449900 488640
rect 340656 488600 449900 488628
rect 340656 488588 340662 488600
rect 449894 488588 449900 488600
rect 449952 488588 449958 488640
rect 105354 488520 105360 488572
rect 105412 488560 105418 488572
rect 215294 488560 215300 488572
rect 105412 488532 215300 488560
rect 105412 488520 105418 488532
rect 215294 488520 215300 488532
rect 215352 488520 215358 488572
rect 220722 488520 220728 488572
rect 220780 488560 220786 488572
rect 330478 488560 330484 488572
rect 220780 488532 330484 488560
rect 220780 488520 220786 488532
rect 330478 488520 330484 488532
rect 330536 488560 330542 488572
rect 440234 488560 440240 488572
rect 330536 488532 440240 488560
rect 330536 488520 330542 488532
rect 440234 488520 440240 488532
rect 440292 488520 440298 488572
rect 79778 488452 79784 488504
rect 79836 488492 79842 488504
rect 92934 488492 92940 488504
rect 79836 488464 92940 488492
rect 79836 488452 79842 488464
rect 92934 488452 92940 488464
rect 92992 488492 92998 488504
rect 188706 488492 188712 488504
rect 92992 488464 188712 488492
rect 92992 488452 92998 488464
rect 188706 488452 188712 488464
rect 188764 488452 188770 488504
rect 231762 488452 231768 488504
rect 231820 488492 231826 488504
rect 340598 488492 340604 488504
rect 231820 488464 340604 488492
rect 231820 488452 231826 488464
rect 340598 488452 340604 488464
rect 340656 488452 340662 488504
rect 407942 488452 407948 488504
rect 408000 488492 408006 488504
rect 423674 488492 423680 488504
rect 408000 488464 423680 488492
rect 408000 488452 408006 488464
rect 423674 488452 423680 488464
rect 423732 488452 423738 488504
rect 79870 488384 79876 488436
rect 79928 488424 79934 488436
rect 94222 488424 94228 488436
rect 79928 488396 94228 488424
rect 79928 488384 79934 488396
rect 94222 488384 94228 488396
rect 94280 488424 94286 488436
rect 188798 488424 188804 488436
rect 94280 488396 188804 488424
rect 94280 488384 94286 488396
rect 188798 488384 188804 488396
rect 188856 488384 188862 488436
rect 408218 488384 408224 488436
rect 408276 488424 408282 488436
rect 422570 488424 422576 488436
rect 408276 488396 422576 488424
rect 408276 488384 408282 488396
rect 422570 488384 422576 488396
rect 422628 488384 422634 488436
rect 79962 488316 79968 488368
rect 80020 488356 80026 488368
rect 95326 488356 95332 488368
rect 80020 488328 95332 488356
rect 80020 488316 80026 488328
rect 95326 488316 95332 488328
rect 95384 488316 95390 488368
rect 312538 488180 312544 488232
rect 312596 488220 312602 488232
rect 408218 488220 408224 488232
rect 312596 488192 408224 488220
rect 312596 488180 312602 488192
rect 408218 488180 408224 488192
rect 408276 488180 408282 488232
rect 318886 488112 318892 488164
rect 318944 488152 318950 488164
rect 427814 488152 427820 488164
rect 318944 488124 427820 488152
rect 318944 488112 318950 488124
rect 427814 488112 427820 488124
rect 427872 488112 427878 488164
rect 188706 488044 188712 488096
rect 188764 488084 188770 488096
rect 202874 488084 202880 488096
rect 188764 488056 202880 488084
rect 188764 488044 188770 488056
rect 202874 488044 202880 488056
rect 202932 488044 202938 488096
rect 326338 488044 326344 488096
rect 326396 488084 326402 488096
rect 434714 488084 434720 488096
rect 326396 488056 434720 488084
rect 326396 488044 326402 488056
rect 434714 488044 434720 488056
rect 434772 488044 434778 488096
rect 188798 487976 188804 488028
rect 188856 488016 188862 488028
rect 204254 488016 204260 488028
rect 188856 487988 204260 488016
rect 188856 487976 188862 487988
rect 204254 487976 204260 487988
rect 204312 487976 204318 488028
rect 360470 487976 360476 488028
rect 360528 488016 360534 488028
rect 470594 488016 470600 488028
rect 360528 487988 470600 488016
rect 360528 487976 360534 487988
rect 470594 487976 470600 487988
rect 470652 487976 470658 488028
rect 102410 487908 102416 487960
rect 102468 487948 102474 487960
rect 211798 487948 211804 487960
rect 102468 487920 211804 487948
rect 102468 487908 102474 487920
rect 211798 487908 211804 487920
rect 211856 487908 211862 487960
rect 219618 487908 219624 487960
rect 219676 487948 219682 487960
rect 281534 487948 281540 487960
rect 219676 487920 281540 487948
rect 219676 487908 219682 487920
rect 281534 487908 281540 487920
rect 281592 487908 281598 487960
rect 345750 487908 345756 487960
rect 345808 487948 345814 487960
rect 455414 487948 455420 487960
rect 345808 487920 455420 487948
rect 345808 487908 345814 487920
rect 455414 487908 455420 487920
rect 455472 487908 455478 487960
rect 135530 487840 135536 487892
rect 135588 487880 135594 487892
rect 244550 487880 244556 487892
rect 135588 487852 244556 487880
rect 135588 487840 135594 487852
rect 244550 487840 244556 487852
rect 244608 487840 244614 487892
rect 355778 487840 355784 487892
rect 355836 487880 355842 487892
rect 465074 487880 465080 487892
rect 355836 487852 465080 487880
rect 355836 487840 355842 487852
rect 465074 487840 465080 487852
rect 465132 487840 465138 487892
rect 125594 487772 125600 487824
rect 125652 487812 125658 487824
rect 235626 487812 235632 487824
rect 125652 487784 235632 487812
rect 125652 487772 125658 487784
rect 235626 487772 235632 487784
rect 235684 487812 235690 487824
rect 235902 487812 235908 487824
rect 235684 487784 235908 487812
rect 235684 487772 235690 487784
rect 235902 487772 235908 487784
rect 235960 487812 235966 487824
rect 235960 487784 238754 487812
rect 235960 487772 235966 487784
rect 97810 487704 97816 487756
rect 97868 487744 97874 487756
rect 207658 487744 207664 487756
rect 97868 487716 207664 487744
rect 97868 487704 97874 487716
rect 207658 487704 207664 487716
rect 207716 487704 207722 487756
rect 105722 487636 105728 487688
rect 105780 487676 105786 487688
rect 215938 487676 215944 487688
rect 105780 487648 215944 487676
rect 105780 487636 105786 487648
rect 215938 487636 215944 487648
rect 215996 487636 216002 487688
rect 104802 487568 104808 487620
rect 104860 487608 104866 487620
rect 214558 487608 214564 487620
rect 104860 487580 214564 487608
rect 104860 487568 104866 487580
rect 214558 487568 214564 487580
rect 214616 487568 214622 487620
rect 99190 487500 99196 487552
rect 99248 487540 99254 487552
rect 209038 487540 209044 487552
rect 99248 487512 209044 487540
rect 99248 487500 99254 487512
rect 209038 487500 209044 487512
rect 209096 487500 209102 487552
rect 100018 487432 100024 487484
rect 100076 487472 100082 487484
rect 210050 487472 210056 487484
rect 100076 487444 210056 487472
rect 100076 487432 100082 487444
rect 210050 487432 210056 487444
rect 210108 487472 210114 487484
rect 211062 487472 211068 487484
rect 210108 487444 211068 487472
rect 210108 487432 210114 487444
rect 211062 487432 211068 487444
rect 211120 487432 211126 487484
rect 238726 487472 238754 487784
rect 241422 487772 241428 487824
rect 241480 487812 241486 487824
rect 350350 487812 350356 487824
rect 241480 487784 350356 487812
rect 241480 487772 241486 487784
rect 350350 487772 350356 487784
rect 350408 487812 350414 487824
rect 459554 487812 459560 487824
rect 350408 487784 459560 487812
rect 350408 487772 350414 487784
rect 459554 487772 459560 487784
rect 459612 487772 459618 487824
rect 318058 487704 318064 487756
rect 318116 487744 318122 487756
rect 426434 487744 426440 487756
rect 318116 487716 426440 487744
rect 318116 487704 318122 487716
rect 426434 487704 426440 487716
rect 426492 487704 426498 487756
rect 320818 487636 320824 487688
rect 320876 487676 320882 487688
rect 430574 487676 430580 487688
rect 320876 487648 430580 487676
rect 320876 487636 320882 487648
rect 430574 487636 430580 487648
rect 430632 487636 430638 487688
rect 320082 487568 320088 487620
rect 320140 487608 320146 487620
rect 429194 487608 429200 487620
rect 320140 487580 429200 487608
rect 320140 487568 320146 487580
rect 429194 487568 429200 487580
rect 429252 487568 429258 487620
rect 322198 487500 322204 487552
rect 322256 487540 322262 487552
rect 432046 487540 432052 487552
rect 322256 487512 432052 487540
rect 322256 487500 322262 487512
rect 432046 487500 432052 487512
rect 432104 487500 432110 487552
rect 345750 487472 345756 487484
rect 238726 487444 345756 487472
rect 345750 487432 345756 487444
rect 345808 487432 345814 487484
rect 103422 487364 103428 487416
rect 103480 487404 103486 487416
rect 213178 487404 213184 487416
rect 103480 487376 213184 487404
rect 103480 487364 103486 487376
rect 213178 487364 213184 487376
rect 213236 487364 213242 487416
rect 250438 487404 250444 487416
rect 238726 487376 250444 487404
rect 101122 487296 101128 487348
rect 101180 487336 101186 487348
rect 211154 487336 211160 487348
rect 101180 487308 211160 487336
rect 101180 487296 101186 487308
rect 211154 487296 211160 487308
rect 211212 487336 211218 487348
rect 212442 487336 212448 487348
rect 211212 487308 212448 487336
rect 211212 487296 211218 487308
rect 212442 487296 212448 487308
rect 212500 487296 212506 487348
rect 140682 487228 140688 487280
rect 140740 487268 140746 487280
rect 238726 487268 238754 487376
rect 250438 487364 250444 487376
rect 250496 487404 250502 487416
rect 251082 487404 251088 487416
rect 250496 487376 251088 487404
rect 250496 487364 250502 487376
rect 251082 487364 251088 487376
rect 251140 487404 251146 487416
rect 360470 487404 360476 487416
rect 251140 487376 360476 487404
rect 251140 487364 251146 487376
rect 360470 487364 360476 487376
rect 360528 487364 360534 487416
rect 244550 487296 244556 487348
rect 244608 487336 244614 487348
rect 245562 487336 245568 487348
rect 244608 487308 245568 487336
rect 244608 487296 244614 487308
rect 245562 487296 245568 487308
rect 245620 487336 245626 487348
rect 355778 487336 355784 487348
rect 245620 487308 355784 487336
rect 245620 487296 245626 487308
rect 355778 487296 355784 487308
rect 355836 487296 355842 487348
rect 140740 487240 238754 487268
rect 140740 487228 140746 487240
rect 323578 487228 323584 487280
rect 323636 487268 323642 487280
rect 433334 487268 433340 487280
rect 323636 487240 433340 487268
rect 323636 487228 323642 487240
rect 433334 487228 433340 487240
rect 433392 487228 433398 487280
rect 130654 487160 130660 487212
rect 130712 487200 130718 487212
rect 241422 487200 241428 487212
rect 130712 487172 241428 487200
rect 130712 487160 130718 487172
rect 241422 487160 241428 487172
rect 241480 487160 241486 487212
rect 324314 487160 324320 487212
rect 324372 487200 324378 487212
rect 324866 487200 324872 487212
rect 324372 487172 324872 487200
rect 324372 487160 324378 487172
rect 324866 487160 324872 487172
rect 324924 487200 324930 487212
rect 434714 487200 434720 487212
rect 324924 487172 434720 487200
rect 324924 487160 324930 487172
rect 434714 487160 434720 487172
rect 434772 487160 434778 487212
rect 212442 486480 212448 486532
rect 212500 486520 212506 486532
rect 247678 486520 247684 486532
rect 212500 486492 247684 486520
rect 212500 486480 212506 486492
rect 247678 486480 247684 486492
rect 247736 486480 247742 486532
rect 187694 486412 187700 486464
rect 187752 486452 187758 486464
rect 241514 486452 241520 486464
rect 187752 486424 241520 486452
rect 187752 486412 187758 486424
rect 241514 486412 241520 486424
rect 241572 486412 241578 486464
rect 244918 486412 244924 486464
rect 244976 486452 244982 486464
rect 318886 486452 318892 486464
rect 244976 486424 318892 486452
rect 244976 486412 244982 486424
rect 318886 486412 318892 486424
rect 318944 486412 318950 486464
rect 187050 485052 187056 485104
rect 187108 485092 187114 485104
rect 261478 485092 261484 485104
rect 187108 485064 261484 485092
rect 187108 485052 187114 485064
rect 261478 485052 261484 485064
rect 261536 485052 261542 485104
rect 261570 485052 261576 485104
rect 261628 485092 261634 485104
rect 297910 485092 297916 485104
rect 261628 485064 297916 485092
rect 261628 485052 261634 485064
rect 297910 485052 297916 485064
rect 297968 485052 297974 485104
rect 211154 484372 211160 484424
rect 211212 484412 211218 484424
rect 580166 484412 580172 484424
rect 211212 484384 580172 484412
rect 211212 484372 211218 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 241514 484304 241520 484356
rect 241572 484344 241578 484356
rect 284938 484344 284944 484356
rect 241572 484316 284944 484344
rect 241572 484304 241578 484316
rect 284938 484304 284944 484316
rect 284996 484304 285002 484356
rect 242802 482332 242808 482384
rect 242860 482372 242866 482384
rect 294690 482372 294696 482384
rect 242860 482344 294696 482372
rect 242860 482332 242866 482344
rect 294690 482332 294696 482344
rect 294748 482332 294754 482384
rect 211062 482264 211068 482316
rect 211120 482304 211126 482316
rect 246114 482304 246120 482316
rect 211120 482276 246120 482304
rect 211120 482264 211126 482276
rect 246114 482264 246120 482276
rect 246172 482264 246178 482316
rect 250346 482264 250352 482316
rect 250404 482304 250410 482316
rect 324314 482304 324320 482316
rect 250404 482276 324320 482304
rect 250404 482264 250410 482276
rect 324314 482264 324320 482276
rect 324372 482264 324378 482316
rect 207658 481040 207664 481092
rect 207716 481080 207722 481092
rect 243538 481080 243544 481092
rect 207716 481052 243544 481080
rect 207716 481040 207722 481052
rect 243538 481040 243544 481052
rect 243596 481040 243602 481092
rect 240134 480972 240140 481024
rect 240192 481012 240198 481024
rect 284110 481012 284116 481024
rect 240192 480984 284116 481012
rect 240192 480972 240198 480984
rect 284110 480972 284116 480984
rect 284168 480972 284174 481024
rect 235994 480904 236000 480956
rect 236052 480944 236058 480956
rect 297450 480944 297456 480956
rect 236052 480916 297456 480944
rect 236052 480904 236058 480916
rect 297450 480904 297456 480916
rect 297508 480904 297514 480956
rect 239950 479544 239956 479596
rect 240008 479584 240014 479596
rect 284018 479584 284024 479596
rect 240008 479556 284024 479584
rect 240008 479544 240014 479556
rect 284018 479544 284024 479556
rect 284076 479544 284082 479596
rect 220722 479476 220728 479528
rect 220780 479516 220786 479528
rect 244274 479516 244280 479528
rect 220780 479488 244280 479516
rect 220780 479476 220786 479488
rect 244274 479476 244280 479488
rect 244332 479476 244338 479528
rect 251634 479476 251640 479528
rect 251692 479516 251698 479528
rect 326338 479516 326344 479528
rect 251692 479488 326344 479516
rect 251692 479476 251698 479488
rect 326338 479476 326344 479488
rect 326396 479476 326402 479528
rect 189074 478796 189080 478848
rect 189132 478836 189138 478848
rect 241882 478836 241888 478848
rect 189132 478808 241888 478836
rect 189132 478796 189138 478808
rect 241882 478796 241888 478808
rect 241940 478796 241946 478848
rect 245838 478796 245844 478848
rect 245896 478836 245902 478848
rect 319438 478836 319444 478848
rect 245896 478808 319444 478836
rect 245896 478796 245902 478808
rect 319438 478796 319444 478808
rect 319496 478796 319502 478848
rect 240042 478184 240048 478236
rect 240100 478224 240106 478236
rect 282362 478224 282368 478236
rect 240100 478196 282368 478224
rect 240100 478184 240106 478196
rect 282362 478184 282368 478196
rect 282420 478184 282426 478236
rect 188246 478116 188252 478168
rect 188304 478156 188310 478168
rect 240870 478156 240876 478168
rect 188304 478128 240876 478156
rect 188304 478116 188310 478128
rect 240870 478116 240876 478128
rect 240928 478116 240934 478168
rect 241882 477980 241888 478032
rect 241940 478020 241946 478032
rect 242802 478020 242808 478032
rect 241940 477992 242808 478020
rect 241940 477980 241946 477992
rect 242802 477980 242808 477992
rect 242860 477980 242866 478032
rect 188614 477436 188620 477488
rect 188672 477476 188678 477488
rect 240134 477476 240140 477488
rect 188672 477448 240140 477476
rect 188672 477436 188678 477448
rect 240134 477436 240140 477448
rect 240192 477436 240198 477488
rect 245562 477436 245568 477488
rect 245620 477476 245626 477488
rect 249794 477476 249800 477488
rect 245620 477448 249800 477476
rect 245620 477436 245626 477448
rect 249794 477436 249800 477448
rect 249852 477436 249858 477488
rect 187602 476756 187608 476808
rect 187660 476796 187666 476808
rect 236362 476796 236368 476808
rect 187660 476768 236368 476796
rect 187660 476756 187666 476768
rect 236362 476756 236368 476768
rect 236420 476756 236426 476808
rect 249150 476756 249156 476808
rect 249208 476796 249214 476808
rect 323578 476796 323584 476808
rect 249208 476768 323584 476796
rect 249208 476756 249214 476768
rect 323578 476756 323584 476768
rect 323636 476756 323642 476808
rect 299106 476416 299112 476468
rect 299164 476456 299170 476468
rect 299382 476456 299388 476468
rect 299164 476428 299388 476456
rect 299164 476416 299170 476428
rect 299382 476416 299388 476428
rect 299440 476416 299446 476468
rect 214558 476008 214564 476060
rect 214616 476048 214622 476060
rect 250346 476048 250352 476060
rect 214616 476020 250352 476048
rect 214616 476008 214622 476020
rect 250346 476008 250352 476020
rect 250404 476008 250410 476060
rect 298646 476008 298652 476060
rect 298704 476048 298710 476060
rect 299198 476048 299204 476060
rect 298704 476020 299204 476048
rect 298704 476008 298710 476020
rect 299198 476008 299204 476020
rect 299256 476048 299262 476060
rect 313918 476048 313924 476060
rect 299256 476020 313924 476048
rect 299256 476008 299262 476020
rect 313918 476008 313924 476020
rect 313976 476008 313982 476060
rect 173250 475464 173256 475516
rect 173308 475504 173314 475516
rect 221090 475504 221096 475516
rect 173308 475476 221096 475504
rect 173308 475464 173314 475476
rect 221090 475464 221096 475476
rect 221148 475464 221154 475516
rect 51810 475396 51816 475448
rect 51868 475436 51874 475448
rect 224126 475436 224132 475448
rect 51868 475408 224132 475436
rect 51868 475396 51874 475408
rect 224126 475396 224132 475408
rect 224184 475396 224190 475448
rect 238110 475396 238116 475448
rect 238168 475436 238174 475448
rect 298646 475436 298652 475448
rect 238168 475408 298652 475436
rect 238168 475396 238174 475408
rect 298646 475396 298652 475408
rect 298704 475396 298710 475448
rect 15838 475328 15844 475380
rect 15896 475368 15902 475380
rect 224034 475368 224040 475380
rect 15896 475340 224040 475368
rect 15896 475328 15902 475340
rect 224034 475328 224040 475340
rect 224092 475328 224098 475380
rect 249058 475328 249064 475380
rect 249116 475368 249122 475380
rect 322198 475368 322204 475380
rect 249116 475340 322204 475368
rect 249116 475328 249122 475340
rect 322198 475328 322204 475340
rect 322256 475328 322262 475380
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 14550 474756 14556 474768
rect 3108 474728 14556 474756
rect 3108 474716 3114 474728
rect 14550 474716 14556 474728
rect 14608 474716 14614 474768
rect 188522 474648 188528 474700
rect 188580 474688 188586 474700
rect 238754 474688 238760 474700
rect 188580 474660 238760 474688
rect 188580 474648 188586 474660
rect 238754 474648 238760 474660
rect 238812 474688 238818 474700
rect 239950 474688 239956 474700
rect 238812 474660 239956 474688
rect 238812 474648 238818 474660
rect 239950 474648 239956 474660
rect 240008 474648 240014 474700
rect 247034 474648 247040 474700
rect 247092 474688 247098 474700
rect 247678 474688 247684 474700
rect 247092 474660 247684 474688
rect 247092 474648 247098 474660
rect 247678 474648 247684 474660
rect 247736 474688 247742 474700
rect 320818 474688 320824 474700
rect 247736 474660 320824 474688
rect 247736 474648 247742 474660
rect 320818 474648 320824 474660
rect 320876 474648 320882 474700
rect 299382 474580 299388 474632
rect 299440 474620 299446 474632
rect 312538 474620 312544 474632
rect 299440 474592 312544 474620
rect 299440 474580 299446 474592
rect 312538 474580 312544 474592
rect 312596 474580 312602 474632
rect 238018 473968 238024 474020
rect 238076 474008 238082 474020
rect 299382 474008 299388 474020
rect 238076 473980 299388 474008
rect 238076 473968 238082 473980
rect 299382 473968 299388 473980
rect 299440 473968 299446 474020
rect 188338 473288 188344 473340
rect 188396 473328 188402 473340
rect 239122 473328 239128 473340
rect 188396 473300 239128 473328
rect 188396 473288 188402 473300
rect 239122 473288 239128 473300
rect 239180 473328 239186 473340
rect 240042 473328 240048 473340
rect 239180 473300 240048 473328
rect 239180 473288 239186 473300
rect 240042 473288 240048 473300
rect 240100 473288 240106 473340
rect 243078 473288 243084 473340
rect 243136 473328 243142 473340
rect 243538 473328 243544 473340
rect 243136 473300 243544 473328
rect 243136 473288 243142 473300
rect 243538 473288 243544 473300
rect 243596 473328 243602 473340
rect 318058 473328 318064 473340
rect 243596 473300 318064 473328
rect 243596 473288 243602 473300
rect 318058 473288 318064 473300
rect 318116 473288 318122 473340
rect 241422 472676 241428 472728
rect 241480 472716 241486 472728
rect 248690 472716 248696 472728
rect 241480 472688 248696 472716
rect 241480 472676 241486 472688
rect 248690 472676 248696 472688
rect 248748 472676 248754 472728
rect 218054 472608 218060 472660
rect 218112 472648 218118 472660
rect 290550 472648 290556 472660
rect 218112 472620 290556 472648
rect 218112 472608 218118 472620
rect 290550 472608 290556 472620
rect 290608 472608 290614 472660
rect 215938 471928 215944 471980
rect 215996 471968 216002 471980
rect 251634 471968 251640 471980
rect 215996 471940 251640 471968
rect 215996 471928 216002 471940
rect 251634 471928 251640 471940
rect 251692 471928 251698 471980
rect 298646 471928 298652 471980
rect 298704 471968 298710 471980
rect 299106 471968 299112 471980
rect 298704 471940 299112 471968
rect 298704 471928 298710 471940
rect 299106 471928 299112 471940
rect 299164 471968 299170 471980
rect 315298 471968 315304 471980
rect 299164 471940 315304 471968
rect 299164 471928 299170 471940
rect 315298 471928 315304 471940
rect 315356 471928 315362 471980
rect 177390 471248 177396 471300
rect 177448 471288 177454 471300
rect 221274 471288 221280 471300
rect 177448 471260 221280 471288
rect 177448 471248 177454 471260
rect 221274 471248 221280 471260
rect 221332 471248 221338 471300
rect 238202 471248 238208 471300
rect 238260 471288 238266 471300
rect 298646 471288 298652 471300
rect 238260 471260 298652 471288
rect 238260 471248 238266 471260
rect 298646 471248 298652 471260
rect 298704 471248 298710 471300
rect 217318 470568 217324 470620
rect 217376 470608 217382 470620
rect 580166 470608 580172 470620
rect 217376 470580 580172 470608
rect 217376 470568 217382 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 216858 469888 216864 469940
rect 216916 469928 216922 469940
rect 392578 469928 392584 469940
rect 216916 469900 392584 469928
rect 216916 469888 216922 469900
rect 392578 469888 392584 469900
rect 392636 469888 392642 469940
rect 216674 469820 216680 469872
rect 216732 469860 216738 469872
rect 402330 469860 402336 469872
rect 216732 469832 402336 469860
rect 216732 469820 216738 469832
rect 402330 469820 402336 469832
rect 402388 469820 402394 469872
rect 186958 469140 186964 469192
rect 187016 469180 187022 469192
rect 261202 469180 261208 469192
rect 187016 469152 261208 469180
rect 187016 469140 187022 469152
rect 261202 469140 261208 469152
rect 261260 469140 261266 469192
rect 261202 468868 261208 468920
rect 261260 468908 261266 468920
rect 261570 468908 261576 468920
rect 261260 468880 261576 468908
rect 261260 468868 261266 468880
rect 261570 468868 261576 468880
rect 261628 468868 261634 468920
rect 213914 468528 213920 468580
rect 213972 468568 213978 468580
rect 523678 468568 523684 468580
rect 213972 468540 523684 468568
rect 213972 468528 213978 468540
rect 523678 468528 523684 468540
rect 523736 468528 523742 468580
rect 215294 468460 215300 468512
rect 215352 468500 215358 468512
rect 533338 468500 533344 468512
rect 215352 468472 533344 468500
rect 215352 468460 215358 468472
rect 533338 468460 533344 468472
rect 533396 468460 533402 468512
rect 218238 467236 218244 467288
rect 218296 467276 218302 467288
rect 298830 467276 298836 467288
rect 218296 467248 298836 467276
rect 218296 467236 218302 467248
rect 298830 467236 298836 467248
rect 298888 467236 298894 467288
rect 77938 467168 77944 467220
rect 77996 467208 78002 467220
rect 236178 467208 236184 467220
rect 77996 467180 236184 467208
rect 77996 467168 78002 467180
rect 236178 467168 236184 467180
rect 236236 467168 236242 467220
rect 214098 467100 214104 467152
rect 214156 467140 214162 467152
rect 580258 467140 580264 467152
rect 214156 467112 580264 467140
rect 214156 467100 214162 467112
rect 580258 467100 580264 467112
rect 580316 467100 580322 467152
rect 218146 465740 218152 465792
rect 218204 465780 218210 465792
rect 397454 465780 397460 465792
rect 218204 465752 397460 465780
rect 218204 465740 218210 465752
rect 397454 465740 397460 465752
rect 397512 465740 397518 465792
rect 215478 465672 215484 465724
rect 215536 465712 215542 465724
rect 527174 465712 527180 465724
rect 215536 465684 527180 465712
rect 215536 465672 215542 465684
rect 527174 465672 527180 465684
rect 527232 465672 527238 465724
rect 218330 464448 218336 464500
rect 218388 464488 218394 464500
rect 409138 464488 409144 464500
rect 218388 464460 409144 464488
rect 218388 464448 218394 464460
rect 409138 464448 409144 464460
rect 409196 464448 409202 464500
rect 214190 464380 214196 464432
rect 214248 464420 214254 464432
rect 503070 464420 503076 464432
rect 214248 464392 503076 464420
rect 214248 464380 214254 464392
rect 503070 464380 503076 464392
rect 503128 464380 503134 464432
rect 212534 464312 212540 464364
rect 212592 464352 212598 464364
rect 515398 464352 515404 464364
rect 212592 464324 515404 464352
rect 212592 464312 212598 464324
rect 515398 464312 515404 464324
rect 515456 464312 515462 464364
rect 51718 463088 51724 463140
rect 51776 463128 51782 463140
rect 222654 463128 222660 463140
rect 51776 463100 222660 463128
rect 51776 463088 51782 463100
rect 222654 463088 222660 463100
rect 222712 463088 222718 463140
rect 236270 463088 236276 463140
rect 236328 463128 236334 463140
rect 408034 463128 408040 463140
rect 236328 463100 408040 463128
rect 236328 463088 236334 463100
rect 408034 463088 408040 463100
rect 408092 463088 408098 463140
rect 216950 463020 216956 463072
rect 217008 463060 217014 463072
rect 402238 463060 402244 463072
rect 217008 463032 402244 463060
rect 217008 463020 217014 463032
rect 402238 463020 402244 463032
rect 402296 463020 402302 463072
rect 212718 462952 212724 463004
rect 212776 462992 212782 463004
rect 549898 462992 549904 463004
rect 212776 462964 549904 462992
rect 212776 462952 212782 462964
rect 549898 462952 549904 462964
rect 549956 462952 549962 463004
rect 3418 462340 3424 462392
rect 3476 462380 3482 462392
rect 226978 462380 226984 462392
rect 3476 462352 226984 462380
rect 3476 462340 3482 462352
rect 226978 462340 226984 462352
rect 227036 462340 227042 462392
rect 217042 461796 217048 461848
rect 217100 461836 217106 461848
rect 393958 461836 393964 461848
rect 217100 461808 393964 461836
rect 217100 461796 217106 461808
rect 393958 461796 393964 461808
rect 394016 461796 394022 461848
rect 3510 461728 3516 461780
rect 3568 461768 3574 461780
rect 225598 461768 225604 461780
rect 3568 461740 225604 461768
rect 3568 461728 3574 461740
rect 225598 461728 225604 461740
rect 225656 461728 225662 461780
rect 215570 461660 215576 461712
rect 215628 461700 215634 461712
rect 505738 461700 505744 461712
rect 215628 461672 505744 461700
rect 215628 461660 215634 461672
rect 505738 461660 505744 461672
rect 505796 461660 505802 461712
rect 216766 461592 216772 461644
rect 216824 461632 216830 461644
rect 542354 461632 542360 461644
rect 216824 461604 542360 461632
rect 216824 461592 216830 461604
rect 542354 461592 542360 461604
rect 542412 461592 542418 461644
rect 215386 460300 215392 460352
rect 215444 460340 215450 460352
rect 502978 460340 502984 460352
rect 215444 460312 502984 460340
rect 215444 460300 215450 460312
rect 502978 460300 502984 460312
rect 503036 460300 503042 460352
rect 214374 460232 214380 460284
rect 214432 460272 214438 460284
rect 503162 460272 503168 460284
rect 214432 460244 503168 460272
rect 214432 460232 214438 460244
rect 503162 460232 503168 460244
rect 503220 460232 503226 460284
rect 212810 460164 212816 460216
rect 212868 460204 212874 460216
rect 519538 460204 519544 460216
rect 212868 460176 519544 460204
rect 212868 460164 212874 460176
rect 519538 460164 519544 460176
rect 519596 460164 519602 460216
rect 213178 459484 213184 459536
rect 213236 459524 213242 459536
rect 248966 459524 248972 459536
rect 213236 459496 248972 459524
rect 213236 459484 213242 459496
rect 248966 459484 248972 459496
rect 249024 459524 249030 459536
rect 249150 459524 249156 459536
rect 249024 459496 249156 459524
rect 249024 459484 249030 459496
rect 249150 459484 249156 459496
rect 249208 459484 249214 459536
rect 204898 459416 204904 459468
rect 204956 459456 204962 459468
rect 238202 459456 238208 459468
rect 204956 459428 238208 459456
rect 204956 459416 204962 459428
rect 238202 459416 238208 459428
rect 238260 459416 238266 459468
rect 205082 459348 205088 459400
rect 205140 459388 205146 459400
rect 238110 459388 238116 459400
rect 205140 459360 238116 459388
rect 205140 459348 205146 459360
rect 238110 459348 238116 459360
rect 238168 459348 238174 459400
rect 237926 458872 237932 458924
rect 237984 458912 237990 458924
rect 238202 458912 238208 458924
rect 237984 458884 238208 458912
rect 237984 458872 237990 458884
rect 238202 458872 238208 458884
rect 238260 458872 238266 458924
rect 246298 458872 246304 458924
rect 246356 458912 246362 458924
rect 371510 458912 371516 458924
rect 246356 458884 371516 458912
rect 246356 458872 246362 458884
rect 371510 458872 371516 458884
rect 371568 458872 371574 458924
rect 260926 458804 260932 458856
rect 260984 458844 260990 458856
rect 309042 458844 309048 458856
rect 260984 458816 309048 458844
rect 260984 458804 260990 458816
rect 309042 458804 309048 458816
rect 309100 458804 309106 458856
rect 298830 458736 298836 458788
rect 298888 458776 298894 458788
rect 329650 458776 329656 458788
rect 298888 458748 329656 458776
rect 298888 458736 298894 458748
rect 329650 458736 329656 458748
rect 329708 458736 329714 458788
rect 295978 458668 295984 458720
rect 296036 458708 296042 458720
rect 346394 458708 346400 458720
rect 296036 458680 346400 458708
rect 296036 458668 296042 458680
rect 346394 458668 346400 458680
rect 346452 458668 346458 458720
rect 298922 458600 298928 458652
rect 298980 458640 298986 458652
rect 354766 458640 354772 458652
rect 298980 458612 354772 458640
rect 298980 458600 298986 458612
rect 354766 458600 354772 458612
rect 354824 458600 354830 458652
rect 299566 458532 299572 458584
rect 299624 458572 299630 458584
rect 359274 458572 359280 458584
rect 299624 458544 359280 458572
rect 299624 458532 299630 458544
rect 359274 458532 359280 458544
rect 359332 458532 359338 458584
rect 260190 458464 260196 458516
rect 260248 458504 260254 458516
rect 321278 458504 321284 458516
rect 260248 458476 321284 458504
rect 260248 458464 260254 458476
rect 321278 458464 321284 458476
rect 321336 458464 321342 458516
rect 297542 458396 297548 458448
rect 297600 458436 297606 458448
rect 363138 458436 363144 458448
rect 297600 458408 363144 458436
rect 297600 458396 297606 458408
rect 363138 458396 363144 458408
rect 363196 458396 363202 458448
rect 299014 458328 299020 458380
rect 299072 458368 299078 458380
rect 367646 458368 367652 458380
rect 299072 458340 367652 458368
rect 299072 458328 299078 458340
rect 367646 458328 367652 458340
rect 367704 458328 367710 458380
rect 237834 458260 237840 458312
rect 237892 458300 237898 458312
rect 238110 458300 238116 458312
rect 237892 458272 238116 458300
rect 237892 458260 237898 458272
rect 238110 458260 238116 458272
rect 238168 458260 238174 458312
rect 254578 458260 254584 458312
rect 254636 458300 254642 458312
rect 379882 458300 379888 458312
rect 254636 458272 379888 458300
rect 254636 458260 254642 458272
rect 379882 458260 379888 458272
rect 379940 458260 379946 458312
rect 14458 457580 14464 457632
rect 14516 457620 14522 457632
rect 227070 457620 227076 457632
rect 14516 457592 227076 457620
rect 14516 457580 14522 457592
rect 227070 457580 227076 457592
rect 227128 457580 227134 457632
rect 3602 457512 3608 457564
rect 3660 457552 3666 457564
rect 224954 457552 224960 457564
rect 3660 457524 224960 457552
rect 3660 457512 3666 457524
rect 224954 457512 224960 457524
rect 225012 457512 225018 457564
rect 213546 457444 213552 457496
rect 213604 457484 213610 457496
rect 501598 457484 501604 457496
rect 213604 457456 501604 457484
rect 213604 457444 213610 457456
rect 501598 457444 501604 457456
rect 501656 457444 501662 457496
rect 241790 457240 241796 457292
rect 241848 457280 241854 457292
rect 312906 457280 312912 457292
rect 241848 457252 312912 457280
rect 241848 457240 241854 457252
rect 312906 457240 312912 457252
rect 312964 457240 312970 457292
rect 232130 457172 232136 457224
rect 232188 457212 232194 457224
rect 325786 457212 325792 457224
rect 232188 457184 325792 457212
rect 232188 457172 232194 457184
rect 325786 457172 325792 457184
rect 325844 457172 325850 457224
rect 243630 457104 243636 457156
rect 243688 457144 243694 457156
rect 338022 457144 338028 457156
rect 243688 457116 338028 457144
rect 243688 457104 243694 457116
rect 338022 457104 338028 457116
rect 338080 457104 338086 457156
rect 242986 457036 242992 457088
rect 243044 457076 243050 457088
rect 342530 457076 342536 457088
rect 243044 457048 342536 457076
rect 243044 457036 243050 457048
rect 342530 457036 342536 457048
rect 342588 457036 342594 457088
rect 232590 456968 232596 457020
rect 232648 457008 232654 457020
rect 334158 457008 334164 457020
rect 232648 456980 334164 457008
rect 232648 456968 232654 456980
rect 334158 456968 334164 456980
rect 334216 456968 334222 457020
rect 241698 456900 241704 456952
rect 241756 456940 241762 456952
rect 350902 456940 350908 456952
rect 241756 456912 350908 456940
rect 241756 456900 241762 456912
rect 350902 456900 350908 456912
rect 350960 456900 350966 456952
rect 231118 456832 231124 456884
rect 231176 456872 231182 456884
rect 376018 456872 376024 456884
rect 231176 456844 376024 456872
rect 231176 456832 231182 456844
rect 376018 456832 376024 456844
rect 376076 456832 376082 456884
rect 211338 456764 211344 456816
rect 211396 456804 211402 456816
rect 580166 456804 580172 456816
rect 211396 456776 580172 456804
rect 211396 456764 211402 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 223206 456220 223212 456272
rect 223264 456260 223270 456272
rect 317414 456260 317420 456272
rect 223264 456232 317420 456260
rect 223264 456220 223270 456232
rect 317414 456220 317420 456232
rect 317472 456220 317478 456272
rect 258074 456152 258080 456204
rect 258132 456192 258138 456204
rect 385310 456192 385316 456204
rect 258132 456164 385316 456192
rect 258132 456152 258138 456164
rect 385310 456152 385316 456164
rect 385368 456152 385374 456204
rect 255774 456084 255780 456136
rect 255832 456124 255838 456136
rect 384114 456124 384120 456136
rect 255832 456096 384120 456124
rect 255832 456084 255838 456096
rect 384114 456084 384120 456096
rect 384172 456084 384178 456136
rect 250070 456016 250076 456068
rect 250128 456056 250134 456068
rect 384206 456056 384212 456068
rect 250128 456028 384212 456056
rect 250128 456016 250134 456028
rect 384206 456016 384212 456028
rect 384264 456016 384270 456068
rect 244734 455948 244740 456000
rect 244792 455988 244798 456000
rect 384022 455988 384028 456000
rect 244792 455960 384028 455988
rect 244792 455948 244798 455960
rect 384022 455948 384028 455960
rect 384080 455948 384086 456000
rect 239030 455880 239036 455932
rect 239088 455920 239094 455932
rect 385034 455920 385040 455932
rect 239088 455892 385040 455920
rect 239088 455880 239094 455892
rect 385034 455880 385040 455892
rect 385092 455880 385098 455932
rect 238938 455812 238944 455864
rect 238996 455852 239002 455864
rect 385402 455852 385408 455864
rect 238996 455824 385408 455852
rect 238996 455812 239002 455824
rect 385402 455812 385408 455824
rect 385460 455812 385466 455864
rect 237558 455744 237564 455796
rect 237616 455784 237622 455796
rect 385218 455784 385224 455796
rect 237616 455756 385224 455784
rect 237616 455744 237622 455756
rect 385218 455744 385224 455756
rect 385276 455744 385282 455796
rect 224954 455676 224960 455728
rect 225012 455716 225018 455728
rect 225414 455716 225420 455728
rect 225012 455688 225420 455716
rect 225012 455676 225018 455688
rect 225414 455676 225420 455688
rect 225472 455716 225478 455728
rect 385494 455716 385500 455728
rect 225472 455688 385500 455716
rect 225472 455676 225478 455688
rect 385494 455676 385500 455688
rect 385552 455676 385558 455728
rect 299658 455608 299664 455660
rect 299716 455648 299722 455660
rect 385126 455648 385132 455660
rect 299716 455620 385132 455648
rect 299716 455608 299722 455620
rect 385126 455608 385132 455620
rect 385184 455608 385190 455660
rect 211522 455540 211528 455592
rect 211580 455580 211586 455592
rect 384298 455580 384304 455592
rect 211580 455552 384304 455580
rect 211580 455540 211586 455552
rect 384298 455540 384304 455552
rect 384356 455540 384362 455592
rect 224034 455472 224040 455524
rect 224092 455512 224098 455524
rect 383562 455512 383568 455524
rect 224092 455484 383568 455512
rect 224092 455472 224098 455484
rect 383562 455472 383568 455484
rect 383620 455472 383626 455524
rect 211430 455404 211436 455456
rect 211488 455444 211494 455456
rect 580258 455444 580264 455456
rect 211488 455416 580264 455444
rect 211488 455404 211494 455416
rect 580258 455404 580264 455416
rect 580316 455404 580322 455456
rect 37918 455336 37924 455388
rect 37976 455376 37982 455388
rect 223758 455376 223764 455388
rect 37976 455348 223764 455376
rect 37976 455336 37982 455348
rect 223758 455336 223764 455348
rect 223816 455376 223822 455388
rect 224034 455376 224040 455388
rect 223816 455348 224040 455376
rect 223816 455336 223822 455348
rect 224034 455336 224040 455348
rect 224092 455336 224098 455388
rect 299842 455336 299848 455388
rect 299900 455376 299906 455388
rect 304166 455376 304172 455388
rect 299900 455348 304172 455376
rect 299900 455336 299906 455348
rect 304166 455336 304172 455348
rect 304224 455336 304230 455388
rect 215662 454792 215668 454844
rect 215720 454832 215726 454844
rect 290458 454832 290464 454844
rect 215720 454804 290464 454832
rect 215720 454792 215726 454804
rect 290458 454792 290464 454804
rect 290516 454792 290522 454844
rect 15930 454724 15936 454776
rect 15988 454764 15994 454776
rect 226610 454764 226616 454776
rect 15988 454736 226616 454764
rect 15988 454724 15994 454736
rect 226610 454724 226616 454736
rect 226668 454724 226674 454776
rect 254486 454724 254492 454776
rect 254544 454764 254550 454776
rect 299842 454764 299848 454776
rect 254544 454736 299848 454764
rect 254544 454724 254550 454736
rect 299842 454724 299848 454736
rect 299900 454724 299906 454776
rect 7558 454656 7564 454708
rect 7616 454696 7622 454708
rect 225506 454696 225512 454708
rect 7616 454668 225512 454696
rect 7616 454656 7622 454668
rect 225506 454656 225512 454668
rect 225564 454656 225570 454708
rect 252554 454656 252560 454708
rect 252612 454696 252618 454708
rect 299566 454696 299572 454708
rect 252612 454668 299572 454696
rect 252612 454656 252618 454668
rect 299566 454656 299572 454668
rect 299624 454656 299630 454708
rect 214006 453500 214012 453552
rect 214064 453540 214070 453552
rect 283558 453540 283564 453552
rect 214064 453512 283564 453540
rect 214064 453500 214070 453512
rect 283558 453500 283564 453512
rect 283616 453500 283622 453552
rect 219526 453432 219532 453484
rect 219584 453472 219590 453484
rect 298738 453472 298744 453484
rect 219584 453444 298744 453472
rect 219584 453432 219590 453444
rect 298738 453432 298744 453444
rect 298796 453432 298802 453484
rect 71774 453364 71780 453416
rect 71832 453404 71838 453416
rect 222286 453404 222292 453416
rect 71832 453376 222292 453404
rect 71832 453364 71838 453376
rect 222286 453364 222292 453376
rect 222344 453364 222350 453416
rect 4798 453296 4804 453348
rect 4856 453336 4862 453348
rect 223574 453336 223580 453348
rect 4856 453308 223580 453336
rect 4856 453296 4862 453308
rect 223574 453296 223580 453308
rect 223632 453296 223638 453348
rect 248598 453296 248604 453348
rect 248656 453336 248662 453348
rect 297542 453336 297548 453348
rect 248656 453308 297548 453336
rect 248656 453296 248662 453308
rect 297542 453296 297548 453308
rect 297600 453296 297606 453348
rect 240778 452548 240784 452600
rect 240836 452588 240842 452600
rect 285030 452588 285036 452600
rect 240836 452560 285036 452588
rect 240836 452548 240842 452560
rect 285030 452548 285036 452560
rect 285088 452548 285094 452600
rect 177298 452072 177304 452124
rect 177356 452112 177362 452124
rect 220998 452112 221004 452124
rect 177356 452084 221004 452112
rect 177356 452072 177362 452084
rect 220998 452072 221004 452084
rect 221056 452072 221062 452124
rect 55858 452004 55864 452056
rect 55916 452044 55922 452056
rect 222378 452044 222384 452056
rect 55916 452016 222384 452044
rect 55916 452004 55922 452016
rect 222378 452004 222384 452016
rect 222436 452004 222442 452056
rect 14550 451936 14556 451988
rect 14608 451976 14614 451988
rect 226886 451976 226892 451988
rect 14608 451948 226892 451976
rect 14608 451936 14614 451948
rect 226886 451936 226892 451948
rect 226944 451936 226950 451988
rect 4982 451868 4988 451920
rect 5040 451908 5046 451920
rect 225138 451908 225144 451920
rect 5040 451880 225144 451908
rect 5040 451868 5046 451880
rect 225138 451868 225144 451880
rect 225196 451868 225202 451920
rect 226242 451868 226248 451920
rect 226300 451908 226306 451920
rect 245746 451908 245752 451920
rect 226300 451880 245752 451908
rect 226300 451868 226306 451880
rect 245746 451868 245752 451880
rect 245804 451868 245810 451920
rect 248046 451868 248052 451920
rect 248104 451908 248110 451920
rect 299750 451908 299756 451920
rect 248104 451880 299756 451908
rect 248104 451868 248110 451880
rect 299750 451868 299756 451880
rect 299808 451868 299814 451920
rect 240318 451256 240324 451308
rect 240376 451296 240382 451308
rect 298002 451296 298008 451308
rect 240376 451268 298008 451296
rect 240376 451256 240382 451268
rect 298002 451256 298008 451268
rect 298060 451256 298066 451308
rect 240870 451188 240876 451240
rect 240928 451228 240934 451240
rect 283650 451228 283656 451240
rect 240928 451200 283656 451228
rect 240928 451188 240934 451200
rect 283650 451188 283656 451200
rect 283708 451188 283714 451240
rect 241698 451052 241704 451104
rect 241756 451092 241762 451104
rect 241974 451092 241980 451104
rect 241756 451064 241980 451092
rect 241756 451052 241762 451064
rect 241974 451052 241980 451064
rect 242032 451052 242038 451104
rect 173158 450712 173164 450764
rect 173216 450752 173222 450764
rect 221090 450752 221096 450764
rect 173216 450724 221096 450752
rect 173216 450712 173222 450724
rect 221090 450712 221096 450724
rect 221148 450712 221154 450764
rect 218698 450644 218704 450696
rect 218756 450684 218762 450696
rect 294598 450684 294604 450696
rect 218756 450656 294604 450684
rect 218756 450644 218762 450656
rect 294598 450644 294604 450656
rect 294656 450644 294662 450696
rect 6178 450576 6184 450628
rect 6236 450616 6242 450628
rect 224770 450616 224776 450628
rect 6236 450588 224776 450616
rect 6236 450576 6242 450588
rect 224770 450576 224776 450588
rect 224828 450576 224834 450628
rect 4890 450508 4896 450560
rect 4948 450548 4954 450560
rect 225322 450548 225328 450560
rect 4948 450520 225328 450548
rect 4948 450508 4954 450520
rect 225322 450508 225328 450520
rect 225380 450508 225386 450560
rect 259822 450508 259828 450560
rect 259880 450548 259886 450560
rect 299014 450548 299020 450560
rect 259880 450520 299020 450548
rect 259880 450508 259886 450520
rect 299014 450508 299020 450520
rect 299072 450508 299078 450560
rect 240686 449896 240692 449948
rect 240744 449936 240750 449948
rect 240870 449936 240876 449948
rect 240744 449908 240876 449936
rect 240744 449896 240750 449908
rect 240870 449896 240876 449908
rect 240928 449896 240934 449948
rect 211798 449828 211804 449880
rect 211856 449868 211862 449880
rect 248506 449868 248512 449880
rect 211856 449840 248512 449868
rect 211856 449828 211862 449840
rect 248506 449828 248512 449840
rect 248564 449828 248570 449880
rect 259546 449828 259552 449880
rect 259604 449868 259610 449880
rect 284478 449868 284484 449880
rect 259604 449840 284484 449868
rect 259604 449828 259610 449840
rect 284478 449828 284484 449840
rect 284536 449828 284542 449880
rect 209038 449760 209044 449812
rect 209096 449800 209102 449812
rect 245010 449800 245016 449812
rect 209096 449772 245016 449800
rect 209096 449760 209102 449772
rect 245010 449760 245016 449772
rect 245068 449760 245074 449812
rect 257890 449760 257896 449812
rect 257948 449800 257954 449812
rect 281994 449800 282000 449812
rect 257948 449772 282000 449800
rect 257948 449760 257954 449772
rect 281994 449760 282000 449772
rect 282052 449760 282058 449812
rect 258626 449692 258632 449744
rect 258684 449732 258690 449744
rect 284294 449732 284300 449744
rect 258684 449704 284300 449732
rect 258684 449692 258690 449704
rect 284294 449692 284300 449704
rect 284352 449692 284358 449744
rect 255682 449624 255688 449676
rect 255740 449664 255746 449676
rect 282178 449664 282184 449676
rect 255740 449636 282184 449664
rect 255740 449624 255746 449636
rect 282178 449624 282184 449636
rect 282236 449624 282242 449676
rect 257338 449556 257344 449608
rect 257396 449596 257402 449608
rect 284846 449596 284852 449608
rect 257396 449568 284852 449596
rect 257396 449556 257402 449568
rect 284846 449556 284852 449568
rect 284904 449556 284910 449608
rect 255130 449488 255136 449540
rect 255188 449528 255194 449540
rect 282270 449528 282276 449540
rect 255188 449500 282276 449528
rect 255188 449488 255194 449500
rect 282270 449488 282276 449500
rect 282328 449488 282334 449540
rect 248506 449420 248512 449472
rect 248564 449460 248570 449472
rect 249058 449460 249064 449472
rect 248564 449432 249064 449460
rect 248564 449420 248570 449432
rect 249058 449420 249064 449432
rect 249116 449420 249122 449472
rect 253474 449420 253480 449472
rect 253532 449460 253538 449472
rect 280982 449460 280988 449472
rect 253532 449432 280988 449460
rect 253532 449420 253538 449432
rect 280982 449420 280988 449432
rect 281040 449420 281046 449472
rect 256234 449352 256240 449404
rect 256292 449392 256298 449404
rect 284386 449392 284392 449404
rect 256292 449364 284392 449392
rect 256292 449352 256298 449364
rect 284386 449352 284392 449364
rect 284444 449352 284450 449404
rect 252370 449284 252376 449336
rect 252428 449324 252434 449336
rect 281810 449324 281816 449336
rect 252428 449296 281816 449324
rect 252428 449284 252434 449296
rect 281810 449284 281816 449296
rect 281868 449284 281874 449336
rect 254302 449216 254308 449268
rect 254360 449256 254366 449268
rect 298922 449256 298928 449268
rect 254360 449228 298928 449256
rect 254360 449216 254366 449228
rect 298922 449216 298928 449228
rect 298980 449216 298986 449268
rect 253750 449148 253756 449200
rect 253808 449188 253814 449200
rect 298830 449188 298836 449200
rect 253808 449160 298836 449188
rect 253808 449148 253814 449160
rect 298830 449148 298836 449160
rect 298888 449148 298894 449200
rect 260650 449080 260656 449132
rect 260708 449120 260714 449132
rect 284570 449120 284576 449132
rect 260708 449092 284576 449120
rect 260708 449080 260714 449092
rect 284570 449080 284576 449092
rect 284628 449080 284634 449132
rect 258994 449012 259000 449064
rect 259052 449052 259058 449064
rect 282086 449052 282092 449064
rect 259052 449024 282092 449052
rect 259052 449012 259058 449024
rect 282086 449012 282092 449024
rect 282144 449012 282150 449064
rect 260098 448944 260104 448996
rect 260156 448984 260162 448996
rect 281902 448984 281908 448996
rect 260156 448956 281908 448984
rect 260156 448944 260162 448956
rect 281902 448944 281908 448956
rect 281960 448944 281966 448996
rect 33778 448468 33784 448520
rect 33836 448508 33842 448520
rect 223206 448508 223212 448520
rect 33836 448480 223212 448508
rect 33836 448468 33842 448480
rect 223206 448468 223212 448480
rect 223264 448468 223270 448520
rect 261478 448468 261484 448520
rect 261536 448508 261542 448520
rect 267090 448508 267096 448520
rect 261536 448480 267096 448508
rect 261536 448468 261542 448480
rect 267090 448468 267096 448480
rect 267148 448508 267154 448520
rect 297358 448508 297364 448520
rect 267148 448480 297364 448508
rect 267148 448468 267154 448480
rect 297358 448468 297364 448480
rect 297416 448468 297422 448520
rect 203518 448400 203524 448452
rect 203576 448440 203582 448452
rect 237466 448440 237472 448452
rect 203576 448412 237472 448440
rect 203576 448400 203582 448412
rect 237466 448400 237472 448412
rect 237524 448440 237530 448452
rect 238018 448440 238024 448452
rect 237524 448412 238024 448440
rect 237524 448400 237530 448412
rect 238018 448400 238024 448412
rect 238076 448400 238082 448452
rect 171778 447856 171784 447908
rect 171836 447896 171842 447908
rect 222562 447896 222568 447908
rect 171836 447868 222568 447896
rect 171836 447856 171842 447868
rect 222562 447856 222568 447868
rect 222620 447856 222626 447908
rect 235902 447856 235908 447908
rect 235960 447896 235966 447908
rect 247954 447896 247960 447908
rect 235960 447868 247960 447896
rect 235960 447856 235966 447868
rect 247954 447856 247960 447868
rect 248012 447856 248018 447908
rect 2866 447788 2872 447840
rect 2924 447828 2930 447840
rect 227254 447828 227260 447840
rect 2924 447800 227260 447828
rect 2924 447788 2930 447800
rect 227254 447788 227260 447800
rect 227312 447788 227318 447840
rect 231762 447788 231768 447840
rect 231820 447828 231826 447840
rect 246850 447828 246856 447840
rect 231820 447800 246856 447828
rect 231820 447788 231826 447800
rect 246850 447788 246856 447800
rect 246908 447788 246914 447840
rect 252094 447788 252100 447840
rect 252152 447828 252158 447840
rect 295978 447828 295984 447840
rect 252152 447800 295984 447828
rect 252152 447788 252158 447800
rect 295978 447788 295984 447800
rect 296036 447788 296042 447840
rect 218054 447312 218060 447364
rect 218112 447352 218118 447364
rect 219066 447352 219072 447364
rect 218112 447324 219072 447352
rect 218112 447312 218118 447324
rect 219066 447312 219072 447324
rect 219124 447312 219130 447364
rect 225414 447312 225420 447364
rect 225472 447352 225478 447364
rect 225690 447352 225696 447364
rect 225472 447324 225696 447352
rect 225472 447312 225478 447324
rect 225690 447312 225696 447324
rect 225748 447312 225754 447364
rect 235994 447312 236000 447364
rect 236052 447352 236058 447364
rect 236454 447352 236460 447364
rect 236052 447324 236460 447352
rect 236052 447312 236058 447324
rect 236454 447312 236460 447324
rect 236512 447312 236518 447364
rect 218238 447244 218244 447296
rect 218296 447284 218302 447296
rect 218790 447284 218796 447296
rect 218296 447256 218796 447284
rect 218296 447244 218302 447256
rect 218790 447244 218796 447256
rect 218848 447244 218854 447296
rect 220998 447244 221004 447296
rect 221056 447284 221062 447296
rect 221826 447284 221832 447296
rect 221056 447256 221832 447284
rect 221056 447244 221062 447256
rect 221826 447244 221832 447256
rect 221884 447244 221890 447296
rect 225138 447244 225144 447296
rect 225196 447284 225202 447296
rect 225966 447284 225972 447296
rect 225196 447256 225972 447284
rect 225196 447244 225202 447256
rect 225966 447244 225972 447256
rect 226024 447244 226030 447296
rect 236270 447244 236276 447296
rect 236328 447284 236334 447296
rect 236730 447284 236736 447296
rect 236328 447256 236736 447284
rect 236328 447244 236334 447256
rect 236730 447244 236736 447256
rect 236788 447244 236794 447296
rect 247678 447108 247684 447160
rect 247736 447148 247742 447160
rect 297358 447148 297364 447160
rect 247736 447120 297364 447148
rect 247736 447108 247742 447120
rect 297358 447108 297364 447120
rect 297416 447108 297422 447160
rect 226702 446836 226708 446888
rect 226760 446876 226766 446888
rect 227070 446876 227076 446888
rect 226760 446848 227076 446876
rect 226760 446836 226766 446848
rect 227070 446836 227076 446848
rect 227128 446876 227134 446888
rect 265894 446876 265900 446888
rect 227128 446848 265900 446876
rect 227128 446836 227134 446848
rect 265894 446836 265900 446848
rect 265952 446836 265958 446888
rect 212626 446768 212632 446820
rect 212684 446808 212690 446820
rect 217318 446808 217324 446820
rect 212684 446780 217324 446808
rect 212684 446768 212690 446780
rect 217318 446768 217324 446780
rect 217376 446768 217382 446820
rect 225046 446768 225052 446820
rect 225104 446808 225110 446820
rect 225598 446808 225604 446820
rect 225104 446780 225604 446808
rect 225104 446768 225110 446780
rect 225598 446768 225604 446780
rect 225656 446808 225662 446820
rect 264698 446808 264704 446820
rect 225656 446780 264704 446808
rect 225656 446768 225662 446780
rect 264698 446768 264704 446780
rect 264756 446768 264762 446820
rect 211154 446700 211160 446752
rect 211212 446740 211218 446752
rect 212350 446740 212356 446752
rect 211212 446712 212356 446740
rect 211212 446700 211218 446712
rect 212350 446700 212356 446712
rect 212408 446700 212414 446752
rect 212534 446700 212540 446752
rect 212592 446740 212598 446752
rect 213178 446740 213184 446752
rect 212592 446712 213184 446740
rect 212592 446700 212598 446712
rect 213178 446700 213184 446712
rect 213236 446700 213242 446752
rect 229462 446700 229468 446752
rect 229520 446740 229526 446752
rect 264514 446740 264520 446752
rect 229520 446712 264520 446740
rect 229520 446700 229526 446712
rect 264514 446700 264520 446712
rect 264572 446700 264578 446752
rect 204898 446632 204904 446684
rect 204956 446672 204962 446684
rect 231394 446672 231400 446684
rect 204956 446644 231400 446672
rect 204956 446632 204962 446644
rect 231394 446632 231400 446644
rect 231452 446632 231458 446684
rect 247126 446632 247132 446684
rect 247184 446672 247190 446684
rect 299198 446672 299204 446684
rect 247184 446644 299204 446672
rect 247184 446632 247190 446644
rect 299198 446632 299204 446644
rect 299256 446632 299262 446684
rect 211430 446564 211436 446616
rect 211488 446604 211494 446616
rect 211798 446604 211804 446616
rect 211488 446576 211804 446604
rect 211488 446564 211494 446576
rect 211798 446564 211804 446576
rect 211856 446564 211862 446616
rect 212810 446564 212816 446616
rect 212868 446604 212874 446616
rect 213454 446604 213460 446616
rect 212868 446576 213460 446604
rect 212868 446564 212874 446576
rect 213454 446564 213460 446576
rect 213512 446564 213518 446616
rect 213914 446564 213920 446616
rect 213972 446604 213978 446616
rect 215110 446604 215116 446616
rect 213972 446576 215116 446604
rect 213972 446564 213978 446576
rect 215110 446564 215116 446576
rect 215168 446564 215174 446616
rect 215570 446564 215576 446616
rect 215628 446604 215634 446616
rect 216214 446604 216220 446616
rect 215628 446576 216220 446604
rect 215628 446564 215634 446576
rect 216214 446564 216220 446576
rect 216272 446564 216278 446616
rect 216674 446564 216680 446616
rect 216732 446604 216738 446616
rect 217318 446604 217324 446616
rect 216732 446576 217324 446604
rect 216732 446564 216738 446576
rect 217318 446564 217324 446576
rect 217376 446564 217382 446616
rect 229002 446564 229008 446616
rect 229060 446604 229066 446616
rect 251726 446604 251732 446616
rect 229060 446576 251732 446604
rect 229060 446564 229066 446576
rect 251726 446564 251732 446576
rect 251784 446564 251790 446616
rect 256786 446564 256792 446616
rect 256844 446604 256850 446616
rect 281718 446604 281724 446616
rect 256844 446576 281724 446604
rect 256844 446564 256850 446576
rect 281718 446564 281724 446576
rect 281776 446564 281782 446616
rect 6178 446496 6184 446548
rect 6236 446536 6242 446548
rect 230842 446536 230848 446548
rect 6236 446508 230848 446536
rect 6236 446496 6242 446508
rect 230842 446496 230848 446508
rect 230900 446496 230906 446548
rect 237926 446496 237932 446548
rect 237984 446536 237990 446548
rect 238570 446536 238576 446548
rect 237984 446508 238576 446536
rect 237984 446496 237990 446508
rect 238570 446496 238576 446508
rect 238628 446496 238634 446548
rect 238938 446496 238944 446548
rect 238996 446536 239002 446548
rect 239950 446536 239956 446548
rect 238996 446508 239956 446536
rect 238996 446496 239002 446508
rect 239950 446496 239956 446508
rect 240008 446496 240014 446548
rect 241514 446496 241520 446548
rect 241572 446536 241578 446548
rect 242434 446536 242440 446548
rect 241572 446508 242440 446536
rect 241572 446496 241578 446508
rect 242434 446496 242440 446508
rect 242492 446496 242498 446548
rect 244366 446496 244372 446548
rect 244424 446536 244430 446548
rect 246298 446536 246304 446548
rect 244424 446508 246304 446536
rect 244424 446496 244430 446508
rect 246298 446496 246304 446508
rect 246356 446496 246362 446548
rect 254394 446496 254400 446548
rect 254452 446536 254458 446548
rect 281626 446536 281632 446548
rect 254452 446508 281632 446536
rect 254452 446496 254458 446508
rect 281626 446496 281632 446508
rect 281684 446496 281690 446548
rect 188982 446428 188988 446480
rect 189040 446468 189046 446480
rect 220630 446468 220636 446480
rect 189040 446440 220636 446468
rect 189040 446428 189046 446440
rect 220630 446428 220636 446440
rect 220688 446428 220694 446480
rect 229094 446428 229100 446480
rect 229152 446468 229158 446480
rect 260834 446468 260840 446480
rect 229152 446440 260840 446468
rect 229152 446428 229158 446440
rect 260834 446428 260840 446440
rect 260892 446428 260898 446480
rect 189994 446360 190000 446412
rect 190052 446400 190058 446412
rect 220906 446400 220912 446412
rect 190052 446372 220912 446400
rect 190052 446360 190058 446372
rect 220906 446360 220912 446372
rect 220964 446360 220970 446412
rect 222562 446360 222568 446412
rect 222620 446400 222626 446412
rect 229646 446400 229652 446412
rect 222620 446372 229652 446400
rect 222620 446360 222626 446372
rect 229646 446360 229652 446372
rect 229704 446360 229710 446412
rect 229738 446360 229744 446412
rect 229796 446400 229802 446412
rect 258442 446400 258448 446412
rect 229796 446372 258448 446400
rect 229796 446360 229802 446372
rect 258442 446360 258448 446372
rect 258500 446360 258506 446412
rect 261754 446360 261760 446412
rect 261812 446400 261818 446412
rect 299842 446400 299848 446412
rect 261812 446372 299848 446400
rect 261812 446360 261818 446372
rect 299842 446360 299848 446372
rect 299900 446360 299906 446412
rect 200850 446292 200856 446344
rect 200908 446332 200914 446344
rect 228358 446332 228364 446344
rect 200908 446304 228364 446332
rect 200908 446292 200914 446304
rect 228358 446292 228364 446304
rect 228416 446292 228422 446344
rect 242894 446292 242900 446344
rect 242952 446332 242958 446344
rect 243538 446332 243544 446344
rect 242952 446304 243544 446332
rect 242952 446292 242958 446304
rect 243538 446292 243544 446304
rect 243596 446292 243602 446344
rect 202414 446224 202420 446276
rect 202472 446264 202478 446276
rect 233050 446264 233056 446276
rect 202472 446236 233056 446264
rect 202472 446224 202478 446236
rect 233050 446224 233056 446236
rect 233108 446224 233114 446276
rect 241606 446224 241612 446276
rect 241664 446264 241670 446276
rect 257430 446264 257436 446276
rect 241664 446236 257436 446264
rect 241664 446224 241670 446236
rect 257430 446224 257436 446236
rect 257488 446224 257494 446276
rect 184198 446156 184204 446208
rect 184256 446196 184262 446208
rect 229186 446196 229192 446208
rect 184256 446168 229192 446196
rect 184256 446156 184262 446168
rect 229186 446156 229192 446168
rect 229244 446156 229250 446208
rect 206554 446088 206560 446140
rect 206612 446128 206618 446140
rect 247494 446128 247500 446140
rect 206612 446100 247500 446128
rect 206612 446088 206618 446100
rect 247494 446088 247500 446100
rect 247552 446088 247558 446140
rect 257614 446088 257620 446140
rect 257672 446128 257678 446140
rect 299382 446128 299388 446140
rect 257672 446100 299388 446128
rect 257672 446088 257678 446100
rect 299382 446088 299388 446100
rect 299440 446088 299446 446140
rect 208210 446020 208216 446072
rect 208268 446060 208274 446072
rect 251818 446060 251824 446072
rect 208268 446032 251824 446060
rect 208268 446020 208274 446032
rect 251818 446020 251824 446032
rect 251876 446020 251882 446072
rect 255406 446020 255412 446072
rect 255464 446060 255470 446072
rect 298646 446060 298652 446072
rect 255464 446032 298652 446060
rect 255464 446020 255470 446032
rect 298646 446020 298652 446032
rect 298704 446020 298710 446072
rect 211246 445952 211252 446004
rect 211304 445992 211310 446004
rect 299290 445992 299296 446004
rect 211304 445964 299296 445992
rect 211304 445952 211310 445964
rect 299290 445952 299296 445964
rect 299348 445952 299354 446004
rect 209866 445884 209872 445936
rect 209924 445924 209930 445936
rect 299014 445924 299020 445936
rect 209924 445896 299020 445924
rect 209924 445884 209930 445896
rect 299014 445884 299020 445896
rect 299072 445884 299078 445936
rect 14458 445816 14464 445868
rect 14516 445856 14522 445868
rect 230014 445856 230020 445868
rect 14516 445828 230020 445856
rect 14516 445816 14522 445828
rect 230014 445816 230020 445828
rect 230072 445816 230078 445868
rect 253198 445816 253204 445868
rect 253256 445856 253262 445868
rect 297358 445856 297364 445868
rect 253256 445828 297364 445856
rect 253256 445816 253262 445828
rect 297358 445816 297364 445828
rect 297416 445816 297422 445868
rect 204162 445748 204168 445800
rect 204220 445788 204226 445800
rect 232222 445788 232228 445800
rect 204220 445760 232228 445788
rect 204220 445748 204226 445760
rect 232222 445748 232228 445760
rect 232280 445748 232286 445800
rect 249886 445748 249892 445800
rect 249944 445788 249950 445800
rect 254578 445788 254584 445800
rect 249944 445760 254584 445788
rect 249944 445748 249950 445760
rect 254578 445748 254584 445760
rect 254636 445748 254642 445800
rect 250070 445544 250076 445596
rect 250128 445584 250134 445596
rect 250990 445584 250996 445596
rect 250128 445556 250996 445584
rect 250128 445544 250134 445556
rect 250990 445544 250996 445556
rect 251048 445544 251054 445596
rect 6270 445408 6276 445460
rect 6328 445448 6334 445460
rect 229462 445448 229468 445460
rect 6328 445420 229468 445448
rect 6328 445408 6334 445420
rect 229462 445408 229468 445420
rect 229520 445408 229526 445460
rect 238754 445408 238760 445460
rect 238812 445448 238818 445460
rect 239674 445448 239680 445460
rect 238812 445420 239680 445448
rect 238812 445408 238818 445420
rect 239674 445408 239680 445420
rect 239732 445408 239738 445460
rect 243078 445408 243084 445460
rect 243136 445448 243142 445460
rect 244090 445448 244096 445460
rect 243136 445420 244096 445448
rect 243136 445408 243142 445420
rect 244090 445408 244096 445420
rect 244148 445408 244154 445460
rect 106918 445340 106924 445392
rect 106976 445380 106982 445392
rect 228542 445380 228548 445392
rect 106976 445352 228548 445380
rect 106976 445340 106982 445352
rect 228542 445340 228548 445352
rect 228600 445340 228606 445392
rect 248966 445340 248972 445392
rect 249024 445380 249030 445392
rect 249610 445380 249616 445392
rect 249024 445352 249616 445380
rect 249024 445340 249030 445352
rect 249610 445340 249616 445352
rect 249668 445340 249674 445392
rect 203610 445272 203616 445324
rect 203668 445312 203674 445324
rect 231118 445312 231124 445324
rect 203668 445284 231124 445312
rect 203668 445272 203674 445284
rect 231118 445272 231124 445284
rect 231176 445272 231182 445324
rect 237558 445272 237564 445324
rect 237616 445312 237622 445324
rect 238294 445312 238300 445324
rect 237616 445284 238300 445312
rect 237616 445272 237622 445284
rect 238294 445272 238300 445284
rect 238352 445272 238358 445324
rect 202322 445204 202328 445256
rect 202380 445244 202386 445256
rect 233602 445244 233608 445256
rect 202380 445216 233608 445244
rect 202380 445204 202386 445216
rect 233602 445204 233608 445216
rect 233660 445204 233666 445256
rect 241790 445204 241796 445256
rect 241848 445244 241854 445256
rect 242710 445244 242716 445256
rect 241848 445216 242716 445244
rect 241848 445204 241854 445216
rect 242710 445204 242716 445216
rect 242768 445204 242774 445256
rect 200758 445136 200764 445188
rect 200816 445176 200822 445188
rect 232590 445176 232596 445188
rect 200816 445148 232596 445176
rect 200816 445136 200822 445148
rect 232590 445136 232596 445148
rect 232648 445176 232654 445188
rect 232774 445176 232780 445188
rect 232648 445148 232780 445176
rect 232648 445136 232654 445148
rect 232774 445136 232780 445148
rect 232832 445136 232838 445188
rect 199378 445068 199384 445120
rect 199436 445108 199442 445120
rect 231946 445108 231952 445120
rect 199436 445080 231952 445108
rect 199436 445068 199442 445080
rect 231946 445068 231952 445080
rect 232004 445068 232010 445120
rect 239398 445068 239404 445120
rect 239456 445108 239462 445120
rect 297634 445108 297640 445120
rect 239456 445080 297640 445108
rect 239456 445068 239462 445080
rect 297634 445068 297640 445080
rect 297692 445068 297698 445120
rect 3694 445000 3700 445052
rect 3752 445040 3758 445052
rect 204898 445040 204904 445052
rect 3752 445012 204904 445040
rect 3752 445000 3758 445012
rect 204898 445000 204904 445012
rect 204956 445000 204962 445052
rect 222378 445000 222384 445052
rect 222436 445040 222442 445052
rect 222930 445040 222936 445052
rect 222436 445012 222936 445040
rect 222436 445000 222442 445012
rect 222930 445000 222936 445012
rect 222988 445000 222994 445052
rect 229646 445000 229652 445052
rect 229704 445040 229710 445052
rect 299474 445040 299480 445052
rect 229704 445012 299480 445040
rect 229704 445000 229710 445012
rect 299474 445000 299480 445012
rect 299532 445000 299538 445052
rect 186958 444932 186964 444984
rect 187016 444972 187022 444984
rect 230290 444972 230296 444984
rect 187016 444944 230296 444972
rect 187016 444932 187022 444944
rect 230290 444932 230296 444944
rect 230348 444932 230354 444984
rect 237190 444932 237196 444984
rect 237248 444972 237254 444984
rect 268286 444972 268292 444984
rect 237248 444944 268292 444972
rect 237248 444932 237254 444944
rect 268286 444932 268292 444944
rect 268344 444932 268350 444984
rect 157978 444864 157984 444916
rect 158036 444904 158042 444916
rect 227806 444904 227812 444916
rect 158036 444876 227812 444904
rect 158036 444864 158042 444876
rect 227806 444864 227812 444876
rect 227864 444864 227870 444916
rect 234430 444864 234436 444916
rect 234488 444904 234494 444916
rect 267366 444904 267372 444916
rect 234488 444876 267372 444904
rect 234488 444864 234494 444876
rect 267366 444864 267372 444876
rect 267424 444864 267430 444916
rect 210142 444796 210148 444848
rect 210200 444836 210206 444848
rect 296530 444836 296536 444848
rect 210200 444808 296536 444836
rect 210200 444796 210206 444808
rect 296530 444796 296536 444808
rect 296588 444796 296594 444848
rect 211338 444728 211344 444780
rect 211396 444768 211402 444780
rect 212074 444768 212080 444780
rect 211396 444740 212080 444768
rect 211396 444728 211402 444740
rect 212074 444728 212080 444740
rect 212132 444728 212138 444780
rect 296438 444768 296444 444780
rect 212184 444740 296444 444768
rect 209314 444660 209320 444712
rect 209372 444700 209378 444712
rect 212184 444700 212212 444740
rect 296438 444728 296444 444740
rect 296496 444728 296502 444780
rect 209372 444672 212212 444700
rect 209372 444660 209378 444672
rect 215478 444660 215484 444712
rect 215536 444700 215542 444712
rect 216490 444700 216496 444712
rect 215536 444672 216496 444700
rect 215536 444660 215542 444672
rect 216490 444660 216496 444672
rect 216548 444660 216554 444712
rect 216582 444660 216588 444712
rect 216640 444700 216646 444712
rect 296346 444700 296352 444712
rect 216640 444672 296352 444700
rect 216640 444660 216646 444672
rect 296346 444660 296352 444672
rect 296404 444660 296410 444712
rect 207658 444592 207664 444644
rect 207716 444632 207722 444644
rect 296254 444632 296260 444644
rect 207716 444604 296260 444632
rect 207716 444592 207722 444604
rect 296254 444592 296260 444604
rect 296312 444592 296318 444644
rect 216858 444524 216864 444576
rect 216916 444564 216922 444576
rect 217594 444564 217600 444576
rect 216916 444536 217600 444564
rect 216916 444524 216922 444536
rect 217594 444524 217600 444536
rect 217652 444524 217658 444576
rect 298830 444564 298836 444576
rect 218026 444536 298836 444564
rect 216950 444456 216956 444508
rect 217008 444496 217014 444508
rect 217870 444496 217876 444508
rect 217008 444468 217876 444496
rect 217008 444456 217014 444468
rect 217870 444456 217876 444468
rect 217928 444456 217934 444508
rect 215294 444388 215300 444440
rect 215352 444428 215358 444440
rect 215938 444428 215944 444440
rect 215352 444400 215944 444428
rect 215352 444388 215358 444400
rect 215938 444388 215944 444400
rect 215996 444388 216002 444440
rect 208762 444320 208768 444372
rect 208820 444360 208826 444372
rect 218026 444360 218054 444536
rect 298830 444524 298836 444536
rect 298888 444524 298894 444576
rect 226978 444456 226984 444508
rect 227036 444496 227042 444508
rect 227530 444496 227536 444508
rect 227036 444468 227536 444496
rect 227036 444456 227042 444468
rect 227530 444456 227536 444468
rect 227588 444496 227594 444508
rect 267274 444496 267280 444508
rect 227588 444468 267280 444496
rect 227588 444456 227594 444468
rect 267274 444456 267280 444468
rect 267332 444456 267338 444508
rect 230290 444388 230296 444440
rect 230348 444428 230354 444440
rect 265986 444428 265992 444440
rect 230348 444400 265992 444428
rect 230348 444388 230354 444400
rect 265986 444388 265992 444400
rect 266044 444388 266050 444440
rect 208820 444332 218054 444360
rect 208820 444320 208826 444332
rect 223666 444320 223672 444372
rect 223724 444320 223730 444372
rect 214190 444116 214196 444168
rect 214248 444156 214254 444168
rect 214834 444156 214840 444168
rect 214248 444128 214840 444156
rect 214248 444116 214254 444128
rect 214834 444116 214840 444128
rect 214892 444116 214898 444168
rect 223684 444100 223712 444320
rect 240318 444252 240324 444304
rect 240376 444292 240382 444304
rect 241054 444292 241060 444304
rect 240376 444264 241060 444292
rect 240376 444252 240382 444264
rect 241054 444252 241060 444264
rect 241112 444252 241118 444304
rect 208486 444048 208492 444100
rect 208544 444088 208550 444100
rect 216582 444088 216588 444100
rect 208544 444060 216588 444088
rect 208544 444048 208550 444060
rect 216582 444048 216588 444060
rect 216640 444048 216646 444100
rect 216674 444048 216680 444100
rect 216732 444088 216738 444100
rect 219434 444088 219440 444100
rect 216732 444060 219440 444088
rect 216732 444048 216738 444060
rect 219434 444048 219440 444060
rect 219492 444048 219498 444100
rect 223666 444048 223672 444100
rect 223724 444048 223730 444100
rect 222470 444020 222476 444032
rect 208366 443992 222476 444020
rect 202230 443844 202236 443896
rect 202288 443884 202294 443896
rect 208366 443884 208394 443992
rect 222470 443980 222476 443992
rect 222528 443980 222534 444032
rect 231486 443952 231492 443964
rect 212460 443924 231492 443952
rect 202288 443856 208394 443884
rect 202288 443844 202294 443856
rect 210326 443844 210332 443896
rect 210384 443884 210390 443896
rect 210878 443884 210884 443896
rect 210384 443856 210884 443884
rect 210384 443844 210390 443856
rect 210878 443844 210884 443856
rect 210936 443844 210942 443896
rect 203518 443776 203524 443828
rect 203576 443816 203582 443828
rect 211154 443816 211160 443828
rect 203576 443788 211160 443816
rect 203576 443776 203582 443788
rect 211154 443776 211160 443788
rect 211212 443776 211218 443828
rect 202598 443708 202604 443760
rect 202656 443748 202662 443760
rect 212460 443748 212488 443924
rect 231486 443912 231492 443924
rect 231544 443912 231550 443964
rect 228726 443884 228732 443896
rect 202656 443720 212488 443748
rect 218026 443856 228732 443884
rect 202656 443708 202662 443720
rect 3602 443640 3608 443692
rect 3660 443680 3666 443692
rect 204162 443680 204168 443692
rect 3660 443652 204168 443680
rect 3660 443640 3666 443652
rect 204162 443640 204168 443652
rect 204220 443640 204226 443692
rect 208118 443640 208124 443692
rect 208176 443680 208182 443692
rect 213086 443680 213092 443692
rect 208176 443652 213092 443680
rect 208176 443640 208182 443652
rect 213086 443640 213092 443652
rect 213144 443640 213150 443692
rect 202046 443572 202052 443624
rect 202104 443612 202110 443624
rect 218026 443612 218054 443856
rect 228726 443844 228732 443856
rect 228784 443844 228790 443896
rect 249150 443844 249156 443896
rect 249208 443884 249214 443896
rect 250806 443884 250812 443896
rect 249208 443856 250812 443884
rect 249208 443844 249214 443856
rect 250806 443844 250812 443856
rect 250864 443844 250870 443896
rect 219158 443776 219164 443828
rect 219216 443816 219222 443828
rect 222746 443816 222752 443828
rect 219216 443788 222752 443816
rect 219216 443776 219222 443788
rect 222746 443776 222752 443788
rect 222804 443776 222810 443828
rect 228450 443776 228456 443828
rect 228508 443816 228514 443828
rect 228508 443788 234614 443816
rect 228508 443776 228514 443788
rect 229554 443748 229560 443760
rect 202104 443584 218054 443612
rect 219268 443720 229560 443748
rect 202104 443572 202110 443584
rect 202782 443504 202788 443556
rect 202840 443544 202846 443556
rect 219268 443544 219296 443720
rect 229554 443708 229560 443720
rect 229612 443708 229618 443760
rect 222746 443640 222752 443692
rect 222804 443680 222810 443692
rect 234246 443680 234252 443692
rect 222804 443652 234252 443680
rect 222804 443640 222810 443652
rect 234246 443640 234252 443652
rect 234304 443640 234310 443692
rect 219342 443572 219348 443624
rect 219400 443612 219406 443624
rect 230474 443612 230480 443624
rect 219400 443584 230480 443612
rect 219400 443572 219406 443584
rect 230474 443572 230480 443584
rect 230532 443572 230538 443624
rect 234586 443612 234614 443788
rect 243170 443776 243176 443828
rect 243228 443816 243234 443828
rect 250898 443816 250904 443828
rect 243228 443788 250904 443816
rect 243228 443776 243234 443788
rect 250898 443776 250904 443788
rect 250956 443776 250962 443828
rect 251082 443776 251088 443828
rect 251140 443816 251146 443828
rect 251726 443816 251732 443828
rect 251140 443788 251732 443816
rect 251140 443776 251146 443788
rect 251726 443776 251732 443788
rect 251784 443776 251790 443828
rect 235902 443708 235908 443760
rect 235960 443748 235966 443760
rect 235960 443720 256694 443748
rect 235960 443708 235966 443720
rect 246758 443640 246764 443692
rect 246816 443680 246822 443692
rect 251082 443680 251088 443692
rect 246816 443652 251088 443680
rect 246816 443640 246822 443652
rect 251082 443640 251088 443652
rect 251140 443640 251146 443692
rect 251174 443640 251180 443692
rect 251232 443680 251238 443692
rect 251232 443652 251956 443680
rect 251232 443640 251238 443652
rect 234586 443584 243584 443612
rect 202840 443516 219296 443544
rect 202840 443504 202846 443516
rect 222470 443504 222476 443556
rect 222528 443544 222534 443556
rect 233970 443544 233976 443556
rect 222528 443516 233976 443544
rect 222528 443504 222534 443516
rect 233970 443504 233976 443516
rect 234028 443504 234034 443556
rect 240410 443504 240416 443556
rect 240468 443544 240474 443556
rect 240468 443516 243308 443544
rect 240468 443504 240474 443516
rect 208366 443448 211108 443476
rect 202874 443300 202880 443352
rect 202932 443340 202938 443352
rect 203886 443340 203892 443352
rect 202932 443312 203892 443340
rect 202932 443300 202938 443312
rect 203886 443300 203892 443312
rect 203944 443300 203950 443352
rect 191098 443232 191104 443284
rect 191156 443272 191162 443284
rect 203426 443272 203432 443284
rect 191156 443244 203432 443272
rect 191156 443232 191162 443244
rect 203426 443232 203432 443244
rect 203484 443232 203490 443284
rect 35158 443028 35164 443080
rect 35216 443068 35222 443080
rect 208366 443068 208394 443448
rect 210326 443368 210332 443420
rect 210384 443368 210390 443420
rect 210786 443408 210792 443420
rect 210712 443380 210792 443408
rect 35216 443040 208394 443068
rect 35216 443028 35222 443040
rect 3418 442960 3424 443012
rect 3476 443000 3482 443012
rect 3476 442972 204254 443000
rect 3476 442960 3482 442972
rect 204226 442728 204254 442972
rect 210344 442728 210372 443368
rect 210712 443068 210740 443380
rect 210786 443368 210792 443380
rect 210844 443368 210850 443420
rect 210878 443368 210884 443420
rect 210936 443368 210942 443420
rect 211080 443408 211108 443448
rect 211154 443436 211160 443488
rect 211212 443476 211218 443488
rect 219158 443476 219164 443488
rect 211212 443448 219164 443476
rect 211212 443436 211218 443448
rect 219158 443436 219164 443448
rect 219216 443436 219222 443488
rect 220446 443436 220452 443488
rect 220504 443476 220510 443488
rect 220504 443448 233832 443476
rect 220504 443436 220510 443448
rect 216674 443408 216680 443420
rect 211080 443380 216680 443408
rect 216674 443368 216680 443380
rect 216732 443368 216738 443420
rect 219434 443368 219440 443420
rect 219492 443408 219498 443420
rect 227898 443408 227904 443420
rect 219492 443380 224954 443408
rect 219492 443368 219498 443380
rect 210896 443272 210924 443368
rect 224926 443340 224954 443380
rect 226306 443380 227904 443408
rect 226306 443340 226334 443380
rect 227898 443368 227904 443380
rect 227956 443368 227962 443420
rect 233694 443368 233700 443420
rect 233752 443368 233758 443420
rect 224926 443312 226334 443340
rect 227686 443312 230474 443340
rect 210896 443244 218054 443272
rect 218026 443136 218054 443244
rect 218026 443108 226334 443136
rect 226306 443068 226334 443108
rect 227686 443068 227714 443312
rect 230446 443204 230474 443312
rect 233712 443272 233740 443368
rect 231826 443244 233740 443272
rect 233804 443272 233832 443448
rect 234586 443448 240824 443476
rect 234586 443272 234614 443448
rect 240410 443408 240416 443420
rect 233804 443244 234614 443272
rect 237346 443380 240416 443408
rect 231826 443204 231854 443244
rect 230446 443176 231854 443204
rect 210712 443040 217824 443068
rect 226306 443040 227714 443068
rect 229940 443040 233234 443068
rect 217796 442864 217824 443040
rect 229940 443000 229968 443040
rect 222166 442972 229968 443000
rect 222166 442932 222194 442972
rect 218026 442904 222194 442932
rect 233206 442932 233234 443040
rect 237346 442932 237374 443380
rect 240410 443368 240416 443380
rect 240468 443368 240474 443420
rect 240686 443368 240692 443420
rect 240744 443368 240750 443420
rect 240704 443000 240732 443368
rect 240796 443204 240824 443448
rect 243170 443408 243176 443420
rect 241486 443380 243176 443408
rect 241486 443204 241514 443380
rect 243170 443368 243176 443380
rect 243228 443368 243234 443420
rect 240796 443176 241514 443204
rect 243280 443204 243308 443516
rect 243446 443436 243452 443488
rect 243504 443436 243510 443488
rect 243464 443272 243492 443436
rect 243556 443408 243584 443584
rect 248874 443572 248880 443624
rect 248932 443612 248938 443624
rect 248932 443584 251404 443612
rect 248932 443572 248938 443584
rect 248966 443504 248972 443556
rect 249024 443544 249030 443556
rect 249024 443516 251312 443544
rect 249024 443504 249030 443516
rect 246206 443436 246212 443488
rect 246264 443476 246270 443488
rect 251174 443476 251180 443488
rect 246264 443448 251180 443476
rect 246264 443436 246270 443448
rect 251174 443436 251180 443448
rect 251232 443436 251238 443488
rect 248874 443408 248880 443420
rect 243556 443380 248880 443408
rect 248874 443368 248880 443380
rect 248932 443368 248938 443420
rect 248966 443368 248972 443420
rect 249024 443368 249030 443420
rect 249150 443368 249156 443420
rect 249208 443368 249214 443420
rect 249518 443368 249524 443420
rect 249576 443408 249582 443420
rect 249576 443380 250760 443408
rect 249576 443368 249582 443380
rect 248984 443272 249012 443368
rect 243464 443244 249012 443272
rect 243280 443176 247034 443204
rect 240704 442972 243768 443000
rect 233206 442904 237374 442932
rect 218026 442864 218054 442904
rect 217796 442836 218054 442864
rect 204226 442700 210372 442728
rect 243740 442592 243768 442972
rect 247006 442932 247034 443176
rect 249168 442932 249196 443368
rect 247006 442904 249196 442932
rect 248386 442632 249794 442660
rect 248386 442592 248414 442632
rect 243740 442564 248414 442592
rect 249766 442456 249794 442632
rect 250732 442524 250760 443380
rect 250806 443368 250812 443420
rect 250864 443368 250870 443420
rect 250898 443368 250904 443420
rect 250956 443368 250962 443420
rect 250824 443136 250852 443368
rect 250916 443204 250944 443368
rect 251284 443272 251312 443516
rect 251376 443340 251404 443584
rect 251928 443476 251956 443652
rect 256666 443544 256694 443720
rect 257430 443640 257436 443692
rect 257488 443680 257494 443692
rect 297542 443680 297548 443692
rect 257488 443652 297548 443680
rect 257488 443640 257494 443652
rect 297542 443640 297548 443652
rect 297600 443640 297606 443692
rect 256970 443572 256976 443624
rect 257028 443612 257034 443624
rect 265250 443612 265256 443624
rect 257028 443584 265256 443612
rect 257028 443572 257034 443584
rect 265250 443572 265256 443584
rect 265308 443572 265314 443624
rect 297450 443544 297456 443556
rect 256666 443516 297456 443544
rect 297450 443504 297456 443516
rect 297508 443504 297514 443556
rect 256970 443476 256976 443488
rect 251928 443448 256976 443476
rect 256970 443436 256976 443448
rect 257028 443436 257034 443488
rect 257246 443436 257252 443488
rect 257304 443476 257310 443488
rect 264606 443476 264612 443488
rect 257304 443448 264612 443476
rect 257304 443436 257310 443448
rect 264606 443436 264612 443448
rect 264664 443436 264670 443488
rect 251726 443368 251732 443420
rect 251784 443408 251790 443420
rect 268470 443408 268476 443420
rect 251784 443380 268476 443408
rect 251784 443368 251790 443380
rect 268470 443368 268476 443380
rect 268528 443368 268534 443420
rect 267182 443340 267188 443352
rect 251376 443312 267188 443340
rect 267182 443300 267188 443312
rect 267240 443300 267246 443352
rect 298554 443272 298560 443284
rect 251284 443244 298560 443272
rect 298554 443232 298560 443244
rect 298612 443232 298618 443284
rect 264330 443204 264336 443216
rect 250916 443176 264336 443204
rect 264330 443164 264336 443176
rect 264388 443164 264394 443216
rect 299106 443136 299112 443148
rect 250824 443108 299112 443136
rect 299106 443096 299112 443108
rect 299164 443096 299170 443148
rect 263870 443028 263876 443080
rect 263928 443068 263934 443080
rect 298002 443068 298008 443080
rect 263928 443040 298008 443068
rect 263928 443028 263934 443040
rect 298002 443028 298008 443040
rect 298060 443028 298066 443080
rect 268378 443000 268384 443012
rect 258046 442972 268384 443000
rect 258046 442524 258074 442972
rect 268378 442960 268384 442972
rect 268436 442960 268442 443012
rect 250732 442496 258074 442524
rect 263870 442456 263876 442468
rect 249766 442428 263876 442456
rect 263870 442416 263876 442428
rect 263928 442416 263934 442468
rect 202966 441464 202972 441516
rect 203024 441504 203030 441516
rect 203702 441504 203708 441516
rect 203024 441476 203708 441504
rect 203024 441464 203030 441476
rect 203702 441464 203708 441476
rect 203760 441464 203766 441516
rect 268378 440172 268384 440224
rect 268436 440212 268442 440224
rect 298002 440212 298008 440224
rect 268436 440184 298008 440212
rect 268436 440172 268442 440184
rect 298002 440172 298008 440184
rect 298060 440172 298066 440224
rect 265250 436024 265256 436076
rect 265308 436064 265314 436076
rect 298002 436064 298008 436076
rect 265308 436036 298008 436064
rect 265308 436024 265314 436036
rect 298002 436024 298008 436036
rect 298060 436024 298066 436076
rect 265986 431876 265992 431928
rect 266044 431916 266050 431928
rect 298002 431916 298008 431928
rect 266044 431888 298008 431916
rect 266044 431876 266050 431888
rect 298002 431876 298008 431888
rect 298060 431876 298066 431928
rect 384298 431876 384304 431928
rect 384356 431916 384362 431928
rect 580166 431916 580172 431928
rect 384356 431888 580172 431916
rect 384356 431876 384362 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 267366 426368 267372 426420
rect 267424 426408 267430 426420
rect 298002 426408 298008 426420
rect 267424 426380 298008 426408
rect 267424 426368 267430 426380
rect 298002 426368 298008 426380
rect 298060 426368 298066 426420
rect 3510 423580 3516 423632
rect 3568 423620 3574 423632
rect 157978 423620 157984 423632
rect 3568 423592 157984 423620
rect 3568 423580 3574 423592
rect 157978 423580 157984 423592
rect 158036 423580 158042 423632
rect 267274 422220 267280 422272
rect 267332 422260 267338 422272
rect 297910 422260 297916 422272
rect 267332 422232 297916 422260
rect 267332 422220 267338 422232
rect 297910 422220 297916 422232
rect 297968 422220 297974 422272
rect 3510 411204 3516 411256
rect 3568 411244 3574 411256
rect 200850 411244 200856 411256
rect 3568 411216 200856 411244
rect 3568 411204 3574 411216
rect 200850 411204 200856 411216
rect 200908 411204 200914 411256
rect 268470 408416 268476 408468
rect 268528 408456 268534 408468
rect 298002 408456 298008 408468
rect 268528 408428 298008 408456
rect 268528 408416 268534 408428
rect 298002 408416 298008 408428
rect 298060 408416 298066 408468
rect 267182 404268 267188 404320
rect 267240 404308 267246 404320
rect 296990 404308 296996 404320
rect 267240 404280 296996 404308
rect 267240 404268 267246 404280
rect 296990 404268 296996 404280
rect 297048 404268 297054 404320
rect 264606 401208 264612 401260
rect 264664 401248 264670 401260
rect 385034 401248 385040 401260
rect 264664 401220 385040 401248
rect 264664 401208 264670 401220
rect 385034 401208 385040 401220
rect 385092 401208 385098 401260
rect 264698 400936 264704 400988
rect 264756 400976 264762 400988
rect 264756 400948 328454 400976
rect 264756 400936 264762 400948
rect 265894 400868 265900 400920
rect 265952 400908 265958 400920
rect 328426 400908 328454 400948
rect 265952 400880 316034 400908
rect 328426 400880 328868 400908
rect 265952 400868 265958 400880
rect 316006 400840 316034 400880
rect 316006 400812 321554 400840
rect 321526 400772 321554 400812
rect 321526 400744 328454 400772
rect 328426 400636 328454 400744
rect 328840 400716 328868 400880
rect 338086 400880 354674 400908
rect 328822 400664 328828 400716
rect 328880 400664 328886 400716
rect 338086 400636 338114 400880
rect 354646 400704 354674 400880
rect 370590 400704 370596 400716
rect 354646 400676 370596 400704
rect 370590 400664 370596 400676
rect 370648 400664 370654 400716
rect 328426 400608 338114 400636
rect 299290 400120 299296 400172
rect 299348 400160 299354 400172
rect 579982 400160 579988 400172
rect 299348 400132 579988 400160
rect 299348 400120 299354 400132
rect 579982 400120 579988 400132
rect 580040 400120 580046 400172
rect 254762 399644 254768 399696
rect 254820 399684 254826 399696
rect 255682 399684 255688 399696
rect 254820 399656 255688 399684
rect 254820 399644 254826 399656
rect 255682 399644 255688 399656
rect 255740 399644 255746 399696
rect 252646 399508 252652 399560
rect 252704 399548 252710 399560
rect 254762 399548 254768 399560
rect 252704 399520 254768 399548
rect 252704 399508 252710 399520
rect 254762 399508 254768 399520
rect 254820 399508 254826 399560
rect 331214 399480 331220 399492
rect 253308 399452 331220 399480
rect 252646 399372 252652 399424
rect 252704 399412 252710 399424
rect 253198 399412 253204 399424
rect 252704 399384 253204 399412
rect 252704 399372 252710 399384
rect 253198 399372 253204 399384
rect 253256 399372 253262 399424
rect 253308 399344 253336 399452
rect 331214 399440 331220 399452
rect 331272 399440 331278 399492
rect 297358 399372 297364 399424
rect 297416 399412 297422 399424
rect 307754 399412 307760 399424
rect 297416 399384 307760 399412
rect 297416 399372 297422 399384
rect 307754 399372 307760 399384
rect 307812 399372 307818 399424
rect 253124 399316 253336 399344
rect 253124 399220 253152 399316
rect 253658 399304 253664 399356
rect 253716 399344 253722 399356
rect 333974 399344 333980 399356
rect 253716 399316 333980 399344
rect 253716 399304 253722 399316
rect 333974 399304 333980 399316
rect 334032 399304 334038 399356
rect 299382 399236 299388 399288
rect 299440 399276 299446 399288
rect 341242 399276 341248 399288
rect 299440 399248 341248 399276
rect 299440 399236 299446 399248
rect 341242 399236 341248 399248
rect 341300 399236 341306 399288
rect 253106 399168 253112 399220
rect 253164 399168 253170 399220
rect 253198 399168 253204 399220
rect 253256 399208 253262 399220
rect 274634 399208 274640 399220
rect 253256 399180 274640 399208
rect 253256 399168 253262 399180
rect 274634 399168 274640 399180
rect 274692 399168 274698 399220
rect 298646 399168 298652 399220
rect 298704 399208 298710 399220
rect 366358 399208 366364 399220
rect 298704 399180 366364 399208
rect 298704 399168 298710 399180
rect 366358 399168 366364 399180
rect 366416 399168 366422 399220
rect 241486 399112 251174 399140
rect 240226 398964 240232 399016
rect 240284 399004 240290 399016
rect 241486 399004 241514 399112
rect 240284 398976 241514 399004
rect 251146 399004 251174 399112
rect 264514 399100 264520 399152
rect 264572 399140 264578 399152
rect 337378 399140 337384 399152
rect 264572 399112 337384 399140
rect 264572 399100 264578 399112
rect 337378 399100 337384 399112
rect 337436 399100 337442 399152
rect 264422 399032 264428 399084
rect 264480 399072 264486 399084
rect 345750 399072 345756 399084
rect 264480 399044 345756 399072
rect 264480 399032 264486 399044
rect 345750 399032 345756 399044
rect 345808 399032 345814 399084
rect 383654 399004 383660 399016
rect 251146 398976 383660 399004
rect 240284 398964 240290 398976
rect 383654 398964 383660 398976
rect 383712 398964 383718 399016
rect 241514 398896 241520 398948
rect 241572 398936 241578 398948
rect 400214 398936 400220 398948
rect 241572 398908 400220 398936
rect 241572 398896 241578 398908
rect 400214 398896 400220 398908
rect 400272 398896 400278 398948
rect 216766 398828 216772 398880
rect 216824 398868 216830 398880
rect 217686 398868 217692 398880
rect 216824 398840 217692 398868
rect 216824 398828 216830 398840
rect 217686 398828 217692 398840
rect 217744 398828 217750 398880
rect 242618 398828 242624 398880
rect 242676 398868 242682 398880
rect 242802 398868 242808 398880
rect 242676 398840 242808 398868
rect 242676 398828 242682 398840
rect 242802 398828 242808 398840
rect 242860 398828 242866 398880
rect 245746 398828 245752 398880
rect 245804 398868 245810 398880
rect 455414 398868 455420 398880
rect 245804 398840 455420 398868
rect 245804 398828 245810 398840
rect 455414 398828 455420 398840
rect 455472 398828 455478 398880
rect 3510 398760 3516 398812
rect 3568 398800 3574 398812
rect 35158 398800 35164 398812
rect 3568 398772 35164 398800
rect 3568 398760 3574 398772
rect 35158 398760 35164 398772
rect 35216 398760 35222 398812
rect 208118 398760 208124 398812
rect 208176 398800 208182 398812
rect 219986 398800 219992 398812
rect 208176 398772 219992 398800
rect 208176 398760 208182 398772
rect 219986 398760 219992 398772
rect 220044 398760 220050 398812
rect 231670 398760 231676 398812
rect 231728 398800 231734 398812
rect 253198 398800 253204 398812
rect 231728 398772 253204 398800
rect 231728 398760 231734 398772
rect 253198 398760 253204 398772
rect 253256 398760 253262 398812
rect 255222 398760 255228 398812
rect 255280 398800 255286 398812
rect 255682 398800 255688 398812
rect 255280 398772 255688 398800
rect 255280 398760 255286 398772
rect 255682 398760 255688 398772
rect 255740 398760 255746 398812
rect 299198 398760 299204 398812
rect 299256 398800 299262 398812
rect 303890 398800 303896 398812
rect 299256 398772 303896 398800
rect 299256 398760 299262 398772
rect 303890 398760 303896 398772
rect 303948 398760 303954 398812
rect 207934 398692 207940 398744
rect 207992 398732 207998 398744
rect 212166 398732 212172 398744
rect 207992 398704 212172 398732
rect 207992 398692 207998 398704
rect 212166 398692 212172 398704
rect 212224 398692 212230 398744
rect 219434 398732 219440 398744
rect 214576 398704 219440 398732
rect 208026 398624 208032 398676
rect 208084 398664 208090 398676
rect 214576 398664 214604 398704
rect 219434 398692 219440 398704
rect 219492 398692 219498 398744
rect 244274 398692 244280 398744
rect 244332 398732 244338 398744
rect 257706 398732 257712 398744
rect 244332 398704 257712 398732
rect 244332 398692 244338 398704
rect 257706 398692 257712 398704
rect 257764 398692 257770 398744
rect 267090 398692 267096 398744
rect 267148 398732 267154 398744
rect 374730 398732 374736 398744
rect 267148 398704 374736 398732
rect 267148 398692 267154 398704
rect 374730 398692 374736 398704
rect 374788 398692 374794 398744
rect 208084 398636 214604 398664
rect 208084 398624 208090 398636
rect 217686 398624 217692 398676
rect 217744 398664 217750 398676
rect 219710 398664 219716 398676
rect 217744 398636 219716 398664
rect 217744 398624 217750 398636
rect 219710 398624 219716 398636
rect 219768 398624 219774 398676
rect 236362 398624 236368 398676
rect 236420 398664 236426 398676
rect 253658 398664 253664 398676
rect 236420 398636 253664 398664
rect 236420 398624 236426 398636
rect 253658 398624 253664 398636
rect 253716 398624 253722 398676
rect 256050 398664 256056 398676
rect 253768 398636 256056 398664
rect 207658 398556 207664 398608
rect 207716 398596 207722 398608
rect 222838 398596 222844 398608
rect 207716 398568 222844 398596
rect 207716 398556 207722 398568
rect 222838 398556 222844 398568
rect 222896 398556 222902 398608
rect 242802 398556 242808 398608
rect 242860 398596 242866 398608
rect 253768 398596 253796 398636
rect 256050 398624 256056 398636
rect 256108 398624 256114 398676
rect 268378 398624 268384 398676
rect 268436 398664 268442 398676
rect 354122 398664 354128 398676
rect 268436 398636 354128 398664
rect 268436 398624 268442 398636
rect 354122 398624 354128 398636
rect 354180 398624 354186 398676
rect 242860 398568 253796 398596
rect 242860 398556 242866 398568
rect 298554 398556 298560 398608
rect 298612 398596 298618 398608
rect 349614 398596 349620 398608
rect 298612 398568 349620 398596
rect 298612 398556 298618 398568
rect 349614 398556 349620 398568
rect 349672 398556 349678 398608
rect 207842 398488 207848 398540
rect 207900 398528 207906 398540
rect 225138 398528 225144 398540
rect 207900 398500 225144 398528
rect 207900 398488 207906 398500
rect 225138 398488 225144 398500
rect 225196 398488 225202 398540
rect 236086 398488 236092 398540
rect 236144 398528 236150 398540
rect 253106 398528 253112 398540
rect 236144 398500 253112 398528
rect 236144 398488 236150 398500
rect 253106 398488 253112 398500
rect 253164 398488 253170 398540
rect 297450 398488 297456 398540
rect 297508 398528 297514 398540
rect 320634 398528 320640 398540
rect 297508 398500 320640 398528
rect 297508 398488 297514 398500
rect 320634 398488 320640 398500
rect 320692 398488 320698 398540
rect 207014 398420 207020 398472
rect 207072 398460 207078 398472
rect 226426 398460 226432 398472
rect 207072 398432 226432 398460
rect 207072 398420 207078 398432
rect 226426 398420 226432 398432
rect 226484 398420 226490 398472
rect 246758 398420 246764 398472
rect 246816 398460 246822 398472
rect 262858 398460 262864 398472
rect 246816 398432 262864 398460
rect 246816 398420 246822 398432
rect 262858 398420 262864 398432
rect 262916 398420 262922 398472
rect 188338 398352 188344 398404
rect 188396 398392 188402 398404
rect 212258 398392 212264 398404
rect 188396 398364 212264 398392
rect 188396 398352 188402 398364
rect 212258 398352 212264 398364
rect 212316 398352 212322 398404
rect 212626 398352 212632 398404
rect 212684 398392 212690 398404
rect 216398 398392 216404 398404
rect 212684 398364 216404 398392
rect 212684 398352 212690 398364
rect 216398 398352 216404 398364
rect 216456 398352 216462 398404
rect 248800 398364 253934 398392
rect 189074 398284 189080 398336
rect 189132 398324 189138 398336
rect 225046 398324 225052 398336
rect 189132 398296 225052 398324
rect 189132 398284 189138 398296
rect 225046 398284 225052 398296
rect 225104 398284 225110 398336
rect 229738 398284 229744 398336
rect 229796 398324 229802 398336
rect 248800 398324 248828 398364
rect 229796 398296 248828 398324
rect 253906 398324 253934 398364
rect 255406 398352 255412 398404
rect 255464 398392 255470 398404
rect 282178 398392 282184 398404
rect 255464 398364 282184 398392
rect 255464 398352 255470 398364
rect 282178 398352 282184 398364
rect 282236 398352 282242 398404
rect 256694 398324 256700 398336
rect 253906 398296 256700 398324
rect 229796 398284 229802 398296
rect 256694 398284 256700 398296
rect 256752 398284 256758 398336
rect 260006 398284 260012 398336
rect 260064 398324 260070 398336
rect 383102 398324 383108 398336
rect 260064 398296 383108 398324
rect 260064 398284 260070 398296
rect 383102 398284 383108 398296
rect 383160 398284 383166 398336
rect 171134 398216 171140 398268
rect 171192 398256 171198 398268
rect 223666 398256 223672 398268
rect 171192 398228 223672 398256
rect 171192 398216 171198 398228
rect 223666 398216 223672 398228
rect 223724 398216 223730 398268
rect 230566 398216 230572 398268
rect 230624 398256 230630 398268
rect 230624 398228 234614 398256
rect 230624 398216 230630 398228
rect 139394 398148 139400 398200
rect 139452 398188 139458 398200
rect 234586 398188 234614 398228
rect 243722 398216 243728 398268
rect 243780 398256 243786 398268
rect 257522 398256 257528 398268
rect 243780 398228 257528 398256
rect 243780 398216 243786 398228
rect 257522 398216 257528 398228
rect 257580 398216 257586 398268
rect 251266 398188 251272 398200
rect 139452 398160 214604 398188
rect 234586 398160 251272 398188
rect 139452 398148 139458 398160
rect 15838 398080 15844 398132
rect 15896 398120 15902 398132
rect 210786 398120 210792 398132
rect 15896 398092 210792 398120
rect 15896 398080 15902 398092
rect 210786 398080 210792 398092
rect 210844 398080 210850 398132
rect 214576 398120 214604 398160
rect 251266 398148 251272 398160
rect 251324 398148 251330 398200
rect 254762 398148 254768 398200
rect 254820 398188 254826 398200
rect 543734 398188 543740 398200
rect 254820 398160 543740 398188
rect 254820 398148 254826 398160
rect 543734 398148 543740 398160
rect 543792 398148 543798 398200
rect 221182 398120 221188 398132
rect 214576 398092 221188 398120
rect 221182 398080 221188 398092
rect 221240 398080 221246 398132
rect 242066 398080 242072 398132
rect 242124 398120 242130 398132
rect 242124 398092 253934 398120
rect 242124 398080 242130 398092
rect 209774 398012 209780 398064
rect 209832 398052 209838 398064
rect 212626 398052 212632 398064
rect 209832 398024 212632 398052
rect 209832 398012 209838 398024
rect 212626 398012 212632 398024
rect 212684 398012 212690 398064
rect 216306 398012 216312 398064
rect 216364 398052 216370 398064
rect 223114 398052 223120 398064
rect 216364 398024 223120 398052
rect 216364 398012 216370 398024
rect 223114 398012 223120 398024
rect 223172 398012 223178 398064
rect 253906 398052 253934 398092
rect 254026 398080 254032 398132
rect 254084 398120 254090 398132
rect 561674 398120 561680 398132
rect 254084 398092 561680 398120
rect 254084 398080 254090 398092
rect 561674 398080 561680 398092
rect 561732 398080 561738 398132
rect 256142 398052 256148 398064
rect 253906 398024 256148 398052
rect 256142 398012 256148 398024
rect 256200 398012 256206 398064
rect 212166 397944 212172 397996
rect 212224 397984 212230 397996
rect 218882 397984 218888 397996
rect 212224 397956 218888 397984
rect 212224 397944 212230 397956
rect 218882 397944 218888 397956
rect 218940 397944 218946 397996
rect 260190 397984 260196 397996
rect 253906 397956 260196 397984
rect 209130 397876 209136 397928
rect 209188 397916 209194 397928
rect 217778 397916 217784 397928
rect 209188 397888 217784 397916
rect 209188 397876 209194 397888
rect 217778 397876 217784 397888
rect 217836 397876 217842 397928
rect 246206 397876 246212 397928
rect 246264 397916 246270 397928
rect 253906 397916 253934 397956
rect 260190 397944 260196 397956
rect 260248 397944 260254 397996
rect 246264 397888 253934 397916
rect 246264 397876 246270 397888
rect 254026 397876 254032 397928
rect 254084 397916 254090 397928
rect 260098 397916 260104 397928
rect 254084 397888 260104 397916
rect 254084 397876 254090 397888
rect 260098 397876 260104 397888
rect 260156 397876 260162 397928
rect 215294 397808 215300 397860
rect 215352 397848 215358 397860
rect 223022 397848 223028 397860
rect 215352 397820 223028 397848
rect 215352 397808 215358 397820
rect 223022 397808 223028 397820
rect 223080 397808 223086 397860
rect 232590 397808 232596 397860
rect 232648 397848 232654 397860
rect 232648 397820 234614 397848
rect 232648 397808 232654 397820
rect 209222 397672 209228 397724
rect 209280 397712 209286 397724
rect 218330 397712 218336 397724
rect 209280 397684 218336 397712
rect 209280 397672 209286 397684
rect 218330 397672 218336 397684
rect 218388 397672 218394 397724
rect 219986 397672 219992 397724
rect 220044 397712 220050 397724
rect 227438 397712 227444 397724
rect 220044 397684 227444 397712
rect 220044 397672 220050 397684
rect 227438 397672 227444 397684
rect 227496 397672 227502 397724
rect 210326 397604 210332 397656
rect 210384 397644 210390 397656
rect 215846 397644 215852 397656
rect 210384 397616 215852 397644
rect 210384 397604 210390 397616
rect 215846 397604 215852 397616
rect 215904 397604 215910 397656
rect 219618 397604 219624 397656
rect 219676 397644 219682 397656
rect 220354 397644 220360 397656
rect 219676 397616 220360 397644
rect 219676 397604 219682 397616
rect 220354 397604 220360 397616
rect 220412 397604 220418 397656
rect 220814 397604 220820 397656
rect 220872 397644 220878 397656
rect 227346 397644 227352 397656
rect 220872 397616 227352 397644
rect 220872 397604 220878 397616
rect 227346 397604 227352 397616
rect 227404 397604 227410 397656
rect 234586 397644 234614 397820
rect 238754 397808 238760 397860
rect 238812 397848 238818 397860
rect 242802 397848 242808 397860
rect 238812 397820 242808 397848
rect 238812 397808 238818 397820
rect 242802 397808 242808 397820
rect 242860 397808 242866 397860
rect 245654 397808 245660 397860
rect 245712 397848 245718 397860
rect 245712 397820 249012 397848
rect 245712 397808 245718 397820
rect 239306 397740 239312 397792
rect 239364 397780 239370 397792
rect 246758 397780 246764 397792
rect 239364 397752 246764 397780
rect 239364 397740 239370 397752
rect 246758 397740 246764 397752
rect 246816 397740 246822 397792
rect 240410 397672 240416 397724
rect 240468 397712 240474 397724
rect 246206 397712 246212 397724
rect 240468 397684 246212 397712
rect 240468 397672 240474 397684
rect 246206 397672 246212 397684
rect 246264 397672 246270 397724
rect 248984 397712 249012 397820
rect 253106 397808 253112 397860
rect 253164 397848 253170 397860
rect 253164 397820 267734 397848
rect 253164 397808 253170 397820
rect 251266 397740 251272 397792
rect 251324 397780 251330 397792
rect 259454 397780 259460 397792
rect 251324 397752 259460 397780
rect 251324 397740 251330 397752
rect 259454 397740 259460 397752
rect 259512 397740 259518 397792
rect 254026 397712 254032 397724
rect 248984 397684 254032 397712
rect 254026 397672 254032 397684
rect 254084 397672 254090 397724
rect 258718 397712 258724 397724
rect 254136 397684 258724 397712
rect 239674 397644 239680 397656
rect 234586 397616 239680 397644
rect 239674 397604 239680 397616
rect 239732 397604 239738 397656
rect 239858 397604 239864 397656
rect 239916 397644 239922 397656
rect 243906 397644 243912 397656
rect 239916 397616 243912 397644
rect 239916 397604 239922 397616
rect 243906 397604 243912 397616
rect 243964 397604 243970 397656
rect 244826 397604 244832 397656
rect 244884 397644 244890 397656
rect 254136 397644 254164 397684
rect 258718 397672 258724 397684
rect 258776 397672 258782 397724
rect 257430 397644 257436 397656
rect 244884 397616 254164 397644
rect 254228 397616 257436 397644
rect 244884 397604 244890 397616
rect 212902 397536 212908 397588
rect 212960 397576 212966 397588
rect 213454 397576 213460 397588
rect 212960 397548 213460 397576
rect 212960 397536 212966 397548
rect 213454 397536 213460 397548
rect 213512 397536 213518 397588
rect 213914 397536 213920 397588
rect 213972 397576 213978 397588
rect 217226 397576 217232 397588
rect 213972 397548 217232 397576
rect 213972 397536 213978 397548
rect 217226 397536 217232 397548
rect 217284 397536 217290 397588
rect 222194 397576 222200 397588
rect 219406 397548 222200 397576
rect 209314 397468 209320 397520
rect 209372 397508 209378 397520
rect 210786 397508 210792 397520
rect 209372 397480 210792 397508
rect 209372 397468 209378 397480
rect 210786 397468 210792 397480
rect 210844 397468 210850 397520
rect 212166 397468 212172 397520
rect 212224 397508 212230 397520
rect 213822 397508 213828 397520
rect 212224 397480 213828 397508
rect 212224 397468 212230 397480
rect 213822 397468 213828 397480
rect 213880 397468 213886 397520
rect 219406 397508 219434 397548
rect 222194 397536 222200 397548
rect 222252 397536 222258 397588
rect 227162 397576 227168 397588
rect 222396 397548 227168 397576
rect 222396 397520 222424 397548
rect 227162 397536 227168 397548
rect 227220 397536 227226 397588
rect 234706 397536 234712 397588
rect 234764 397576 234770 397588
rect 240042 397576 240048 397588
rect 234764 397548 240048 397576
rect 234764 397536 234770 397548
rect 240042 397536 240048 397548
rect 240100 397536 240106 397588
rect 240962 397536 240968 397588
rect 241020 397576 241026 397588
rect 246942 397576 246948 397588
rect 241020 397548 246948 397576
rect 241020 397536 241026 397548
rect 246942 397536 246948 397548
rect 247000 397536 247006 397588
rect 216692 397480 219434 397508
rect 212902 397400 212908 397452
rect 212960 397440 212966 397452
rect 216692 397440 216720 397480
rect 220354 397468 220360 397520
rect 220412 397508 220418 397520
rect 220906 397508 220912 397520
rect 220412 397480 220912 397508
rect 220412 397468 220418 397480
rect 220906 397468 220912 397480
rect 220964 397468 220970 397520
rect 222378 397468 222384 397520
rect 222436 397468 222442 397520
rect 226426 397468 226432 397520
rect 226484 397508 226490 397520
rect 227806 397508 227812 397520
rect 226484 397480 227812 397508
rect 226484 397468 226490 397480
rect 227806 397468 227812 397480
rect 227864 397468 227870 397520
rect 238202 397468 238208 397520
rect 238260 397508 238266 397520
rect 242526 397508 242532 397520
rect 238260 397480 242532 397508
rect 238260 397468 238266 397480
rect 242526 397468 242532 397480
rect 242584 397468 242590 397520
rect 243170 397468 243176 397520
rect 243228 397508 243234 397520
rect 254228 397508 254256 397616
rect 257430 397604 257436 397616
rect 257488 397604 257494 397656
rect 267706 397644 267734 397820
rect 525794 397644 525800 397656
rect 267706 397616 525800 397644
rect 525794 397604 525800 397616
rect 525852 397604 525858 397656
rect 254302 397536 254308 397588
rect 254360 397576 254366 397588
rect 564434 397576 564440 397588
rect 254360 397548 564440 397576
rect 254360 397536 254366 397548
rect 564434 397536 564440 397548
rect 564492 397536 564498 397588
rect 243228 397480 254256 397508
rect 243228 397468 243234 397480
rect 256786 397468 256792 397520
rect 256844 397508 256850 397520
rect 582374 397508 582380 397520
rect 256844 397480 582380 397508
rect 256844 397468 256850 397480
rect 582374 397468 582380 397480
rect 582432 397468 582438 397520
rect 212960 397412 216720 397440
rect 212960 397400 212966 397412
rect 237466 397400 237472 397452
rect 237524 397440 237530 397452
rect 238386 397440 238392 397452
rect 237524 397412 238392 397440
rect 237524 397400 237530 397412
rect 238386 397400 238392 397412
rect 238444 397400 238450 397452
rect 210786 397332 210792 397384
rect 210844 397372 210850 397384
rect 224678 397372 224684 397384
rect 210844 397344 224684 397372
rect 210844 397332 210850 397344
rect 224678 397332 224684 397344
rect 224736 397332 224742 397384
rect 37274 397264 37280 397316
rect 37332 397304 37338 397316
rect 213270 397304 213276 397316
rect 37332 397276 213276 397304
rect 37332 397264 37338 397276
rect 213270 397264 213276 397276
rect 213328 397264 213334 397316
rect 245930 397264 245936 397316
rect 245988 397304 245994 397316
rect 257338 397304 257344 397316
rect 245988 397276 257344 397304
rect 245988 397264 245994 397276
rect 257338 397264 257344 397276
rect 257396 397264 257402 397316
rect 212534 397196 212540 397248
rect 212592 397236 212598 397248
rect 213362 397236 213368 397248
rect 212592 397208 213368 397236
rect 212592 397196 212598 397208
rect 213362 397196 213368 397208
rect 213420 397196 213426 397248
rect 198734 397128 198740 397180
rect 198792 397168 198798 397180
rect 225782 397168 225788 397180
rect 198792 397140 225788 397168
rect 198792 397128 198798 397140
rect 225782 397128 225788 397140
rect 225840 397128 225846 397180
rect 234246 397128 234252 397180
rect 234304 397168 234310 397180
rect 234304 397140 234614 397168
rect 234304 397128 234310 397140
rect 162854 397060 162860 397112
rect 162912 397100 162918 397112
rect 215294 397100 215300 397112
rect 162912 397072 215300 397100
rect 162912 397060 162918 397072
rect 215294 397060 215300 397072
rect 215352 397060 215358 397112
rect 151814 396992 151820 397044
rect 151872 397032 151878 397044
rect 212902 397032 212908 397044
rect 151872 397004 212908 397032
rect 151872 396992 151878 397004
rect 212902 396992 212908 397004
rect 212960 396992 212966 397044
rect 212994 396992 213000 397044
rect 213052 397032 213058 397044
rect 213362 397032 213368 397044
rect 213052 397004 213368 397032
rect 213052 396992 213058 397004
rect 213362 396992 213368 397004
rect 213420 396992 213426 397044
rect 214098 396992 214104 397044
rect 214156 397032 214162 397044
rect 214558 397032 214564 397044
rect 214156 397004 214564 397032
rect 214156 396992 214162 397004
rect 214558 396992 214564 397004
rect 214616 396992 214622 397044
rect 218054 396992 218060 397044
rect 218112 397032 218118 397044
rect 218882 397032 218888 397044
rect 218112 397004 218888 397032
rect 218112 396992 218118 397004
rect 218882 396992 218888 397004
rect 218940 396992 218946 397044
rect 144914 396924 144920 396976
rect 144972 396964 144978 396976
rect 221642 396964 221648 396976
rect 144972 396936 221648 396964
rect 144972 396924 144978 396936
rect 221642 396924 221648 396936
rect 221700 396924 221706 396976
rect 131114 396856 131120 396908
rect 131172 396896 131178 396908
rect 131172 396868 214880 396896
rect 131172 396856 131178 396868
rect 40034 396788 40040 396840
rect 40092 396828 40098 396840
rect 212534 396828 212540 396840
rect 40092 396800 212540 396828
rect 40092 396788 40098 396800
rect 212534 396788 212540 396800
rect 212592 396788 212598 396840
rect 210142 396720 210148 396772
rect 210200 396760 210206 396772
rect 210602 396760 210608 396772
rect 210200 396732 210608 396760
rect 210200 396720 210206 396732
rect 210602 396720 210608 396732
rect 210660 396720 210666 396772
rect 211246 396720 211252 396772
rect 211304 396760 211310 396772
rect 211982 396760 211988 396772
rect 211304 396732 211988 396760
rect 211304 396720 211310 396732
rect 211982 396720 211988 396732
rect 212040 396720 212046 396772
rect 212718 396720 212724 396772
rect 212776 396760 212782 396772
rect 213730 396760 213736 396772
rect 212776 396732 213736 396760
rect 212776 396720 212782 396732
rect 213730 396720 213736 396732
rect 213788 396720 213794 396772
rect 209866 396652 209872 396704
rect 209924 396692 209930 396704
rect 210418 396692 210424 396704
rect 209924 396664 210424 396692
rect 209924 396652 209930 396664
rect 210418 396652 210424 396664
rect 210476 396652 210482 396704
rect 211614 396652 211620 396704
rect 211672 396692 211678 396704
rect 211890 396692 211896 396704
rect 211672 396664 211896 396692
rect 211672 396652 211678 396664
rect 211890 396652 211896 396664
rect 211948 396652 211954 396704
rect 212994 396652 213000 396704
rect 213052 396692 213058 396704
rect 213638 396692 213644 396704
rect 213052 396664 213644 396692
rect 213052 396652 213058 396664
rect 213638 396652 213644 396664
rect 213696 396652 213702 396704
rect 214852 396692 214880 396868
rect 218146 396856 218152 396908
rect 218204 396896 218210 396908
rect 218790 396896 218796 396908
rect 218204 396868 218796 396896
rect 218204 396856 218210 396868
rect 218790 396856 218796 396868
rect 218848 396856 218854 396908
rect 219434 396856 219440 396908
rect 219492 396896 219498 396908
rect 220078 396896 220084 396908
rect 219492 396868 220084 396896
rect 219492 396856 219498 396868
rect 220078 396856 220084 396868
rect 220136 396856 220142 396908
rect 222378 396856 222384 396908
rect 222436 396896 222442 396908
rect 222654 396896 222660 396908
rect 222436 396868 222660 396896
rect 222436 396856 222442 396868
rect 222654 396856 222660 396868
rect 222712 396856 222718 396908
rect 234586 396896 234614 397140
rect 237374 397128 237380 397180
rect 237432 397168 237438 397180
rect 237926 397168 237932 397180
rect 237432 397140 237932 397168
rect 237432 397128 237438 397140
rect 237926 397128 237932 397140
rect 237984 397128 237990 397180
rect 237650 396992 237656 397044
rect 237708 397032 237714 397044
rect 237926 397032 237932 397044
rect 237708 397004 237932 397032
rect 237708 396992 237714 397004
rect 237926 396992 237932 397004
rect 237984 396992 237990 397044
rect 307754 396896 307760 396908
rect 234586 396868 307760 396896
rect 307754 396856 307760 396868
rect 307812 396856 307818 396908
rect 215294 396788 215300 396840
rect 215352 396828 215358 396840
rect 215352 396800 218744 396828
rect 215352 396788 215358 396800
rect 215478 396720 215484 396772
rect 215536 396760 215542 396772
rect 215938 396760 215944 396772
rect 215536 396732 215944 396760
rect 215536 396720 215542 396732
rect 215938 396720 215944 396732
rect 215996 396720 216002 396772
rect 218422 396720 218428 396772
rect 218480 396760 218486 396772
rect 218606 396760 218612 396772
rect 218480 396732 218612 396760
rect 218480 396720 218486 396732
rect 218606 396720 218612 396732
rect 218664 396720 218670 396772
rect 218716 396760 218744 396800
rect 219710 396788 219716 396840
rect 219768 396828 219774 396840
rect 220170 396828 220176 396840
rect 219768 396800 220176 396828
rect 219768 396788 219774 396800
rect 220170 396788 220176 396800
rect 220228 396788 220234 396840
rect 222562 396788 222568 396840
rect 222620 396828 222626 396840
rect 222838 396828 222844 396840
rect 222620 396800 222844 396828
rect 222620 396788 222626 396800
rect 222838 396788 222844 396800
rect 222896 396788 222902 396840
rect 223850 396788 223856 396840
rect 223908 396828 223914 396840
rect 224310 396828 224316 396840
rect 223908 396800 224316 396828
rect 223908 396788 223914 396800
rect 224310 396788 224316 396800
rect 224368 396788 224374 396840
rect 236730 396788 236736 396840
rect 236788 396828 236794 396840
rect 339494 396828 339500 396840
rect 236788 396800 339500 396828
rect 236788 396788 236794 396800
rect 339494 396788 339500 396800
rect 339552 396788 339558 396840
rect 223390 396760 223396 396772
rect 218716 396732 223396 396760
rect 223390 396720 223396 396732
rect 223448 396720 223454 396772
rect 241146 396720 241152 396772
rect 241204 396760 241210 396772
rect 396074 396760 396080 396772
rect 241204 396732 396080 396760
rect 241204 396720 241210 396732
rect 396074 396720 396080 396732
rect 396132 396720 396138 396772
rect 220538 396692 220544 396704
rect 214852 396664 220544 396692
rect 220538 396652 220544 396664
rect 220596 396652 220602 396704
rect 221090 396652 221096 396704
rect 221148 396692 221154 396704
rect 221550 396692 221556 396704
rect 221148 396664 221556 396692
rect 221148 396652 221154 396664
rect 221550 396652 221556 396664
rect 221608 396652 221614 396704
rect 224310 396652 224316 396704
rect 224368 396692 224374 396704
rect 224770 396692 224776 396704
rect 224368 396664 224776 396692
rect 224368 396652 224374 396664
rect 224770 396652 224776 396664
rect 224828 396652 224834 396704
rect 210510 396624 210516 396636
rect 209976 396596 210516 396624
rect 209976 396568 210004 396596
rect 210510 396584 210516 396596
rect 210568 396584 210574 396636
rect 211338 396584 211344 396636
rect 211396 396624 211402 396636
rect 212074 396624 212080 396636
rect 211396 396596 212080 396624
rect 211396 396584 211402 396596
rect 212074 396584 212080 396596
rect 212132 396584 212138 396636
rect 212902 396584 212908 396636
rect 212960 396624 212966 396636
rect 213546 396624 213552 396636
rect 212960 396596 213552 396624
rect 212960 396584 212966 396596
rect 213546 396584 213552 396596
rect 213604 396584 213610 396636
rect 214190 396584 214196 396636
rect 214248 396624 214254 396636
rect 215110 396624 215116 396636
rect 214248 396596 215116 396624
rect 214248 396584 214254 396596
rect 215110 396584 215116 396596
rect 215168 396584 215174 396636
rect 215754 396584 215760 396636
rect 215812 396624 215818 396636
rect 216490 396624 216496 396636
rect 215812 396596 216496 396624
rect 215812 396584 215818 396596
rect 216490 396584 216496 396596
rect 216548 396584 216554 396636
rect 218238 396584 218244 396636
rect 218296 396624 218302 396636
rect 219250 396624 219256 396636
rect 218296 396596 219256 396624
rect 218296 396584 218302 396596
rect 219250 396584 219256 396596
rect 219308 396584 219314 396636
rect 219802 396584 219808 396636
rect 219860 396624 219866 396636
rect 220446 396624 220452 396636
rect 219860 396596 220452 396624
rect 219860 396584 219866 396596
rect 220446 396584 220452 396596
rect 220504 396584 220510 396636
rect 220998 396584 221004 396636
rect 221056 396624 221062 396636
rect 221826 396624 221832 396636
rect 221056 396596 221832 396624
rect 221056 396584 221062 396596
rect 221826 396584 221832 396596
rect 221884 396584 221890 396636
rect 223758 396584 223764 396636
rect 223816 396624 223822 396636
rect 224862 396624 224868 396636
rect 223816 396596 224868 396624
rect 223816 396584 223822 396596
rect 224862 396584 224868 396596
rect 224920 396584 224926 396636
rect 232498 396584 232504 396636
rect 232556 396624 232562 396636
rect 232556 396596 232728 396624
rect 232556 396584 232562 396596
rect 209958 396516 209964 396568
rect 210016 396516 210022 396568
rect 210050 396516 210056 396568
rect 210108 396556 210114 396568
rect 210970 396556 210976 396568
rect 210108 396528 210976 396556
rect 210108 396516 210114 396528
rect 210970 396516 210976 396528
rect 211028 396516 211034 396568
rect 211430 396516 211436 396568
rect 211488 396556 211494 396568
rect 212442 396556 212448 396568
rect 211488 396528 212448 396556
rect 211488 396516 211494 396528
rect 212442 396516 212448 396528
rect 212500 396516 212506 396568
rect 214374 396516 214380 396568
rect 214432 396556 214438 396568
rect 215202 396556 215208 396568
rect 214432 396528 215208 396556
rect 214432 396516 214438 396528
rect 215202 396516 215208 396528
rect 215260 396516 215266 396568
rect 215570 396516 215576 396568
rect 215628 396556 215634 396568
rect 216582 396556 216588 396568
rect 215628 396528 216588 396556
rect 215628 396516 215634 396528
rect 216582 396516 216588 396528
rect 216640 396516 216646 396568
rect 216858 396516 216864 396568
rect 216916 396556 216922 396568
rect 217870 396556 217876 396568
rect 216916 396528 217876 396556
rect 216916 396516 216922 396528
rect 217870 396516 217876 396528
rect 217928 396516 217934 396568
rect 218330 396516 218336 396568
rect 218388 396556 218394 396568
rect 218790 396556 218796 396568
rect 218388 396528 218796 396556
rect 218388 396516 218394 396528
rect 218790 396516 218796 396528
rect 218848 396516 218854 396568
rect 219618 396516 219624 396568
rect 219676 396556 219682 396568
rect 220630 396556 220636 396568
rect 219676 396528 220636 396556
rect 219676 396516 219682 396528
rect 220630 396516 220636 396528
rect 220688 396516 220694 396568
rect 221274 396516 221280 396568
rect 221332 396556 221338 396568
rect 221918 396556 221924 396568
rect 221332 396528 221924 396556
rect 221332 396516 221338 396528
rect 221918 396516 221924 396528
rect 221976 396516 221982 396568
rect 222470 396516 222476 396568
rect 222528 396556 222534 396568
rect 223298 396556 223304 396568
rect 222528 396528 223304 396556
rect 222528 396516 222534 396528
rect 223298 396516 223304 396528
rect 223356 396516 223362 396568
rect 224034 396516 224040 396568
rect 224092 396556 224098 396568
rect 224402 396556 224408 396568
rect 224092 396528 224408 396556
rect 224092 396516 224098 396528
rect 224402 396516 224408 396528
rect 224460 396516 224466 396568
rect 232700 396500 232728 396596
rect 242158 396584 242164 396636
rect 242216 396624 242222 396636
rect 242216 396596 242296 396624
rect 242216 396584 242222 396596
rect 213914 396448 213920 396500
rect 213972 396488 213978 396500
rect 215018 396488 215024 396500
rect 213972 396460 215024 396488
rect 213972 396448 213978 396460
rect 215018 396448 215024 396460
rect 215076 396448 215082 396500
rect 218698 396448 218704 396500
rect 218756 396488 218762 396500
rect 219158 396488 219164 396500
rect 218756 396460 219164 396488
rect 218756 396448 218762 396460
rect 219158 396448 219164 396460
rect 219216 396448 219222 396500
rect 219894 396448 219900 396500
rect 219952 396488 219958 396500
rect 220262 396488 220268 396500
rect 219952 396460 220268 396488
rect 219952 396448 219958 396460
rect 220262 396448 220268 396460
rect 220320 396448 220326 396500
rect 221366 396448 221372 396500
rect 221424 396488 221430 396500
rect 222102 396488 222108 396500
rect 221424 396460 222108 396488
rect 221424 396448 221430 396460
rect 222102 396448 222108 396460
rect 222160 396448 222166 396500
rect 232682 396448 232688 396500
rect 232740 396448 232746 396500
rect 209774 396380 209780 396432
rect 209832 396420 209838 396432
rect 210602 396420 210608 396432
rect 209832 396392 210608 396420
rect 209832 396380 209838 396392
rect 210602 396380 210608 396392
rect 210660 396380 210666 396432
rect 213178 396380 213184 396432
rect 213236 396420 213242 396432
rect 215294 396420 215300 396432
rect 213236 396392 215300 396420
rect 213236 396380 213242 396392
rect 215294 396380 215300 396392
rect 215352 396380 215358 396432
rect 217042 396380 217048 396432
rect 217100 396420 217106 396432
rect 217594 396420 217600 396432
rect 217100 396392 217600 396420
rect 217100 396380 217106 396392
rect 217594 396380 217600 396392
rect 217652 396380 217658 396432
rect 218514 396380 218520 396432
rect 218572 396420 218578 396432
rect 219066 396420 219072 396432
rect 218572 396392 219072 396420
rect 218572 396380 218578 396392
rect 219066 396380 219072 396392
rect 219124 396380 219130 396432
rect 242268 396420 242296 396596
rect 242342 396420 242348 396432
rect 242268 396392 242348 396420
rect 242342 396380 242348 396392
rect 242400 396380 242406 396432
rect 215662 396312 215668 396364
rect 215720 396352 215726 396364
rect 216122 396352 216128 396364
rect 215720 396324 216128 396352
rect 215720 396312 215726 396324
rect 216122 396312 216128 396324
rect 216180 396312 216186 396364
rect 217226 396312 217232 396364
rect 217284 396352 217290 396364
rect 217962 396352 217968 396364
rect 217284 396324 217968 396352
rect 217284 396312 217290 396324
rect 217962 396312 217968 396324
rect 218020 396312 218026 396364
rect 218330 396312 218336 396364
rect 218388 396352 218394 396364
rect 218974 396352 218980 396364
rect 218388 396324 218980 396352
rect 218388 396312 218394 396324
rect 218974 396312 218980 396324
rect 219032 396312 219038 396364
rect 217134 396244 217140 396296
rect 217192 396284 217198 396296
rect 217410 396284 217416 396296
rect 217192 396256 217416 396284
rect 217192 396244 217198 396256
rect 217410 396244 217416 396256
rect 217468 396244 217474 396296
rect 219986 396176 219992 396228
rect 220044 396216 220050 396228
rect 220722 396216 220728 396228
rect 220044 396188 220728 396216
rect 220044 396176 220050 396188
rect 220722 396176 220728 396188
rect 220780 396176 220786 396228
rect 220906 396176 220912 396228
rect 220964 396216 220970 396228
rect 222010 396216 222016 396228
rect 220964 396188 222016 396216
rect 220964 396176 220970 396188
rect 222010 396176 222016 396188
rect 222068 396176 222074 396228
rect 244182 396108 244188 396160
rect 244240 396148 244246 396160
rect 245378 396148 245384 396160
rect 244240 396120 245384 396148
rect 244240 396108 244246 396120
rect 245378 396108 245384 396120
rect 245436 396108 245442 396160
rect 210418 396040 210424 396092
rect 210476 396080 210482 396092
rect 210786 396080 210792 396092
rect 210476 396052 210792 396080
rect 210476 396040 210482 396052
rect 210786 396040 210792 396052
rect 210844 396040 210850 396092
rect 210234 395972 210240 396024
rect 210292 396012 210298 396024
rect 211062 396012 211068 396024
rect 210292 395984 211068 396012
rect 210292 395972 210298 395984
rect 211062 395972 211068 395984
rect 211120 395972 211126 396024
rect 217318 395972 217324 396024
rect 217376 396012 217382 396024
rect 217686 396012 217692 396024
rect 217376 395984 217692 396012
rect 217376 395972 217382 395984
rect 217686 395972 217692 395984
rect 217744 395972 217750 396024
rect 220078 395972 220084 396024
rect 220136 396012 220142 396024
rect 226886 396012 226892 396024
rect 220136 395984 226892 396012
rect 220136 395972 220142 395984
rect 226886 395972 226892 395984
rect 226944 395972 226950 396024
rect 204898 395836 204904 395888
rect 204956 395876 204962 395888
rect 224126 395876 224132 395888
rect 204956 395848 224132 395876
rect 204956 395836 204962 395848
rect 224126 395836 224132 395848
rect 224184 395836 224190 395888
rect 230842 395836 230848 395888
rect 230900 395876 230906 395888
rect 231486 395876 231492 395888
rect 230900 395848 231492 395876
rect 230900 395836 230906 395848
rect 231486 395836 231492 395848
rect 231544 395836 231550 395888
rect 218054 395808 218060 395820
rect 209976 395780 218060 395808
rect 115934 395564 115940 395616
rect 115992 395604 115998 395616
rect 209976 395604 210004 395780
rect 218054 395768 218060 395780
rect 218112 395768 218118 395820
rect 231946 395768 231952 395820
rect 232004 395808 232010 395820
rect 232866 395808 232872 395820
rect 232004 395780 232872 395808
rect 232004 395768 232010 395780
rect 232866 395768 232872 395780
rect 232924 395768 232930 395820
rect 218146 395740 218152 395752
rect 115992 395576 210004 395604
rect 210160 395712 218152 395740
rect 115992 395564 115998 395576
rect 109034 395496 109040 395548
rect 109092 395536 109098 395548
rect 210160 395536 210188 395712
rect 218146 395700 218152 395712
rect 218204 395700 218210 395752
rect 246758 395700 246764 395752
rect 246816 395740 246822 395752
rect 372614 395740 372620 395752
rect 246816 395712 372620 395740
rect 246816 395700 246822 395712
rect 372614 395700 372620 395712
rect 372672 395700 372678 395752
rect 215938 395632 215944 395684
rect 215996 395672 216002 395684
rect 216306 395672 216312 395684
rect 215996 395644 216312 395672
rect 215996 395632 216002 395644
rect 216306 395632 216312 395644
rect 216364 395632 216370 395684
rect 247678 395632 247684 395684
rect 247736 395672 247742 395684
rect 248046 395672 248052 395684
rect 247736 395644 248052 395672
rect 247736 395632 247742 395644
rect 248046 395632 248052 395644
rect 248104 395632 248110 395684
rect 249242 395632 249248 395684
rect 249300 395672 249306 395684
rect 499574 395672 499580 395684
rect 249300 395644 499580 395672
rect 249300 395632 249306 395644
rect 499574 395632 499580 395644
rect 499632 395632 499638 395684
rect 214466 395564 214472 395616
rect 214524 395604 214530 395616
rect 214650 395604 214656 395616
rect 214524 395576 214656 395604
rect 214524 395564 214530 395576
rect 214650 395564 214656 395576
rect 214708 395564 214714 395616
rect 250346 395564 250352 395616
rect 250404 395604 250410 395616
rect 514754 395604 514760 395616
rect 250404 395576 514760 395604
rect 250404 395564 250410 395576
rect 514754 395564 514760 395576
rect 514812 395564 514818 395616
rect 216674 395536 216680 395548
rect 109092 395508 210188 395536
rect 210344 395508 216680 395536
rect 109092 395496 109098 395508
rect 93854 395428 93860 395480
rect 93912 395468 93918 395480
rect 210344 395468 210372 395508
rect 216674 395496 216680 395508
rect 216732 395496 216738 395548
rect 251450 395496 251456 395548
rect 251508 395536 251514 395548
rect 528554 395536 528560 395548
rect 251508 395508 528560 395536
rect 251508 395496 251514 395508
rect 528554 395496 528560 395508
rect 528612 395496 528618 395548
rect 93912 395440 210372 395468
rect 93912 395428 93918 395440
rect 214466 395428 214472 395480
rect 214524 395468 214530 395480
rect 214926 395468 214932 395480
rect 214524 395440 214932 395468
rect 214524 395428 214530 395440
rect 214926 395428 214932 395440
rect 214984 395428 214990 395480
rect 252002 395428 252008 395480
rect 252060 395468 252066 395480
rect 535454 395468 535460 395480
rect 252060 395440 535460 395468
rect 252060 395428 252066 395440
rect 535454 395428 535460 395440
rect 535512 395428 535518 395480
rect 86954 395360 86960 395412
rect 87012 395400 87018 395412
rect 214742 395400 214748 395412
rect 87012 395372 214748 395400
rect 87012 395360 87018 395372
rect 214742 395360 214748 395372
rect 214800 395360 214806 395412
rect 253198 395360 253204 395412
rect 253256 395400 253262 395412
rect 549254 395400 549260 395412
rect 253256 395372 549260 395400
rect 253256 395360 253262 395372
rect 549254 395360 549260 395372
rect 549312 395360 549318 395412
rect 77294 395292 77300 395344
rect 77352 395332 77358 395344
rect 216398 395332 216404 395344
rect 77352 395304 216404 395332
rect 77352 395292 77358 395304
rect 216398 395292 216404 395304
rect 216456 395292 216462 395344
rect 255222 395292 255228 395344
rect 255280 395332 255286 395344
rect 571334 395332 571340 395344
rect 255280 395304 571340 395332
rect 255280 395292 255286 395304
rect 571334 395292 571340 395304
rect 571392 395292 571398 395344
rect 240318 395088 240324 395140
rect 240376 395128 240382 395140
rect 240962 395128 240968 395140
rect 240376 395100 240968 395128
rect 240376 395088 240382 395100
rect 240962 395088 240968 395100
rect 241020 395088 241026 395140
rect 242986 395088 242992 395140
rect 243044 395128 243050 395140
rect 243722 395128 243728 395140
rect 243044 395100 243728 395128
rect 243044 395088 243050 395100
rect 243722 395088 243728 395100
rect 243780 395088 243786 395140
rect 248690 395020 248696 395072
rect 248748 395060 248754 395072
rect 249242 395060 249248 395072
rect 248748 395032 249248 395060
rect 248748 395020 248754 395032
rect 249242 395020 249248 395032
rect 249300 395020 249306 395072
rect 214006 394952 214012 395004
rect 214064 394992 214070 395004
rect 214834 394992 214840 395004
rect 214064 394964 214840 394992
rect 214064 394952 214070 394964
rect 214834 394952 214840 394964
rect 214892 394952 214898 395004
rect 213270 394884 213276 394936
rect 213328 394924 213334 394936
rect 213822 394924 213828 394936
rect 213328 394896 213828 394924
rect 213328 394884 213334 394896
rect 213822 394884 213828 394896
rect 213880 394884 213886 394936
rect 253934 394748 253940 394800
rect 253992 394788 253998 394800
rect 254762 394788 254768 394800
rect 253992 394760 254768 394788
rect 253992 394748 253998 394760
rect 254762 394748 254768 394760
rect 254820 394748 254826 394800
rect 235994 394612 236000 394664
rect 236052 394652 236058 394664
rect 244182 394652 244188 394664
rect 236052 394624 244188 394652
rect 236052 394612 236058 394624
rect 244182 394612 244188 394624
rect 244240 394612 244246 394664
rect 244550 394612 244556 394664
rect 244608 394652 244614 394664
rect 244826 394652 244832 394664
rect 244608 394624 244832 394652
rect 244608 394612 244614 394624
rect 244826 394612 244832 394624
rect 244884 394612 244890 394664
rect 247034 394612 247040 394664
rect 247092 394652 247098 394664
rect 247092 394624 250392 394652
rect 247092 394612 247098 394624
rect 236822 394544 236828 394596
rect 236880 394584 236886 394596
rect 244090 394584 244096 394596
rect 236880 394556 244096 394584
rect 236880 394544 236886 394556
rect 244090 394544 244096 394556
rect 244148 394544 244154 394596
rect 244366 394544 244372 394596
rect 244424 394584 244430 394596
rect 244918 394584 244924 394596
rect 244424 394556 244924 394584
rect 244424 394544 244430 394556
rect 244918 394544 244924 394556
rect 244976 394544 244982 394596
rect 249886 394544 249892 394596
rect 249944 394584 249950 394596
rect 250254 394584 250260 394596
rect 249944 394556 250260 394584
rect 249944 394544 249950 394556
rect 250254 394544 250260 394556
rect 250312 394544 250318 394596
rect 250364 394584 250392 394624
rect 251542 394612 251548 394664
rect 251600 394652 251606 394664
rect 252186 394652 252192 394664
rect 251600 394624 252192 394652
rect 251600 394612 251606 394624
rect 252186 394612 252192 394624
rect 252244 394612 252250 394664
rect 253934 394612 253940 394664
rect 253992 394652 253998 394664
rect 254578 394652 254584 394664
rect 253992 394624 254584 394652
rect 253992 394612 253998 394624
rect 254578 394612 254584 394624
rect 254636 394612 254642 394664
rect 255958 394584 255964 394596
rect 250364 394556 255964 394584
rect 255958 394544 255964 394556
rect 256016 394544 256022 394596
rect 237466 394476 237472 394528
rect 237524 394516 237530 394528
rect 243998 394516 244004 394528
rect 237524 394488 244004 394516
rect 237524 394476 237530 394488
rect 243998 394476 244004 394488
rect 244056 394476 244062 394528
rect 244274 394476 244280 394528
rect 244332 394516 244338 394528
rect 244642 394516 244648 394528
rect 244332 394488 244648 394516
rect 244332 394476 244338 394488
rect 244642 394476 244648 394488
rect 244700 394476 244706 394528
rect 245746 394476 245752 394528
rect 245804 394516 245810 394528
rect 246022 394516 246028 394528
rect 245804 394488 246028 394516
rect 245804 394476 245810 394488
rect 246022 394476 246028 394488
rect 246080 394476 246086 394528
rect 250162 394476 250168 394528
rect 250220 394516 250226 394528
rect 250806 394516 250812 394528
rect 250220 394488 250812 394516
rect 250220 394476 250226 394488
rect 250806 394476 250812 394488
rect 250864 394476 250870 394528
rect 251542 394476 251548 394528
rect 251600 394516 251606 394528
rect 251910 394516 251916 394528
rect 251600 394488 251916 394516
rect 251600 394476 251606 394488
rect 251910 394476 251916 394488
rect 251968 394476 251974 394528
rect 252830 394476 252836 394528
rect 252888 394516 252894 394528
rect 253198 394516 253204 394528
rect 252888 394488 253204 394516
rect 252888 394476 252894 394488
rect 253198 394476 253204 394488
rect 253256 394476 253262 394528
rect 254118 394476 254124 394528
rect 254176 394516 254182 394528
rect 254394 394516 254400 394528
rect 254176 394488 254400 394516
rect 254176 394476 254182 394488
rect 254394 394476 254400 394488
rect 254452 394476 254458 394528
rect 227254 394408 227260 394460
rect 227312 394408 227318 394460
rect 234338 394408 234344 394460
rect 234396 394448 234402 394460
rect 307846 394448 307852 394460
rect 234396 394420 307852 394448
rect 234396 394408 234402 394420
rect 307846 394408 307852 394420
rect 307904 394408 307910 394460
rect 209038 394204 209044 394256
rect 209096 394244 209102 394256
rect 219434 394244 219440 394256
rect 209096 394216 219440 394244
rect 209096 394204 209102 394216
rect 219434 394204 219440 394216
rect 219492 394204 219498 394256
rect 225598 394244 225604 394256
rect 222488 394216 225604 394244
rect 195974 394136 195980 394188
rect 196032 394176 196038 394188
rect 222488 394176 222516 394216
rect 225598 394204 225604 394216
rect 225656 394204 225662 394256
rect 227272 394244 227300 394408
rect 235166 394340 235172 394392
rect 235224 394380 235230 394392
rect 318794 394380 318800 394392
rect 235224 394352 235396 394380
rect 235224 394340 235230 394352
rect 228450 394272 228456 394324
rect 228508 394312 228514 394324
rect 228726 394312 228732 394324
rect 228508 394284 228732 394312
rect 228508 394272 228514 394284
rect 228726 394272 228732 394284
rect 228784 394272 228790 394324
rect 233786 394272 233792 394324
rect 233844 394312 233850 394324
rect 234062 394312 234068 394324
rect 233844 394284 234068 394312
rect 233844 394272 233850 394284
rect 234062 394272 234068 394284
rect 234120 394272 234126 394324
rect 234706 394272 234712 394324
rect 234764 394312 234770 394324
rect 235258 394312 235264 394324
rect 234764 394284 235264 394312
rect 234764 394272 234770 394284
rect 235258 394272 235264 394284
rect 235316 394272 235322 394324
rect 227346 394244 227352 394256
rect 227272 394216 227352 394244
rect 227346 394204 227352 394216
rect 227404 394204 227410 394256
rect 235368 394244 235396 394352
rect 243924 394352 318800 394380
rect 240134 394272 240140 394324
rect 240192 394312 240198 394324
rect 241146 394312 241152 394324
rect 240192 394284 241152 394312
rect 240192 394272 240198 394284
rect 241146 394272 241152 394284
rect 241204 394272 241210 394324
rect 241514 394272 241520 394324
rect 241572 394312 241578 394324
rect 241790 394312 241796 394324
rect 241572 394284 241796 394312
rect 241572 394272 241578 394284
rect 241790 394272 241796 394284
rect 241848 394272 241854 394324
rect 242894 394272 242900 394324
rect 242952 394312 242958 394324
rect 243170 394312 243176 394324
rect 242952 394284 243176 394312
rect 242952 394272 242958 394284
rect 243170 394272 243176 394284
rect 243228 394272 243234 394324
rect 235368 394216 242296 394244
rect 196032 394148 222516 394176
rect 196032 394136 196038 394148
rect 224126 394136 224132 394188
rect 224184 394176 224190 394188
rect 224494 394176 224500 394188
rect 224184 394148 224500 394176
rect 224184 394136 224190 394148
rect 224494 394136 224500 394148
rect 224552 394136 224558 394188
rect 231946 394136 231952 394188
rect 232004 394176 232010 394188
rect 232222 394176 232228 394188
rect 232004 394148 232228 394176
rect 232004 394136 232010 394148
rect 232222 394136 232228 394148
rect 232280 394136 232286 394188
rect 234614 394136 234620 394188
rect 234672 394176 234678 394188
rect 235166 394176 235172 394188
rect 234672 394148 235172 394176
rect 234672 394136 234678 394148
rect 235166 394136 235172 394148
rect 235224 394136 235230 394188
rect 239030 394136 239036 394188
rect 239088 394176 239094 394188
rect 239088 394148 240272 394176
rect 239088 394136 239094 394148
rect 168374 394068 168380 394120
rect 168432 394108 168438 394120
rect 223482 394108 223488 394120
rect 168432 394080 223488 394108
rect 168432 394068 168438 394080
rect 223482 394068 223488 394080
rect 223540 394068 223546 394120
rect 232406 394068 232412 394120
rect 232464 394108 232470 394120
rect 232590 394108 232596 394120
rect 232464 394080 232596 394108
rect 232464 394068 232470 394080
rect 232590 394068 232596 394080
rect 232648 394068 232654 394120
rect 234982 394068 234988 394120
rect 235040 394108 235046 394120
rect 235350 394108 235356 394120
rect 235040 394080 235356 394108
rect 235040 394068 235046 394080
rect 235350 394068 235356 394080
rect 235408 394068 235414 394120
rect 240244 394108 240272 394148
rect 241698 394136 241704 394188
rect 241756 394176 241762 394188
rect 242158 394176 242164 394188
rect 241756 394148 242164 394176
rect 241756 394136 241762 394148
rect 242158 394136 242164 394148
rect 242216 394136 242222 394188
rect 242268 394176 242296 394216
rect 242802 394204 242808 394256
rect 242860 394244 242866 394256
rect 243538 394244 243544 394256
rect 242860 394216 243544 394244
rect 242860 394204 242866 394216
rect 243538 394204 243544 394216
rect 243596 394204 243602 394256
rect 243924 394176 243952 394352
rect 318794 394340 318800 394352
rect 318852 394340 318858 394392
rect 244182 394272 244188 394324
rect 244240 394312 244246 394324
rect 329834 394312 329840 394324
rect 244240 394284 329840 394312
rect 244240 394272 244246 394284
rect 329834 394272 329840 394284
rect 329892 394272 329898 394324
rect 244090 394204 244096 394256
rect 244148 394244 244154 394256
rect 340874 394244 340880 394256
rect 244148 394216 340880 394244
rect 244148 394204 244154 394216
rect 340874 394204 340880 394216
rect 340932 394204 340938 394256
rect 242268 394148 243952 394176
rect 243998 394136 244004 394188
rect 244056 394176 244062 394188
rect 347774 394176 347780 394188
rect 244056 394148 347780 394176
rect 244056 394136 244062 394148
rect 347774 394136 347780 394148
rect 347832 394136 347838 394188
rect 240244 394080 242388 394108
rect 143534 394000 143540 394052
rect 143592 394040 143598 394052
rect 221458 394040 221464 394052
rect 143592 394012 221464 394040
rect 143592 394000 143598 394012
rect 221458 394000 221464 394012
rect 221516 394000 221522 394052
rect 228542 394000 228548 394052
rect 228600 394040 228606 394052
rect 234614 394040 234620 394052
rect 228600 394012 234620 394040
rect 228600 394000 228606 394012
rect 234614 394000 234620 394012
rect 234672 394000 234678 394052
rect 235994 394000 236000 394052
rect 236052 394040 236058 394052
rect 236914 394040 236920 394052
rect 236052 394012 236920 394040
rect 236052 394000 236058 394012
rect 236914 394000 236920 394012
rect 236972 394000 236978 394052
rect 241974 394000 241980 394052
rect 242032 394040 242038 394052
rect 242250 394040 242256 394052
rect 242032 394012 242256 394040
rect 242032 394000 242038 394012
rect 242250 394000 242256 394012
rect 242308 394000 242314 394052
rect 242360 394040 242388 394080
rect 242710 394068 242716 394120
rect 242768 394108 242774 394120
rect 365714 394108 365720 394120
rect 242768 394080 365720 394108
rect 242768 394068 242774 394080
rect 365714 394068 365720 394080
rect 365772 394068 365778 394120
rect 368474 394040 368480 394052
rect 242360 394012 368480 394040
rect 368474 394000 368480 394012
rect 368532 394000 368538 394052
rect 63494 393932 63500 393984
rect 63552 393972 63558 393984
rect 212442 393972 212448 393984
rect 63552 393944 212448 393972
rect 63552 393932 63558 393944
rect 212442 393932 212448 393944
rect 212500 393932 212506 393984
rect 219434 393932 219440 393984
rect 219492 393972 219498 393984
rect 220170 393972 220176 393984
rect 219492 393944 220176 393972
rect 219492 393932 219498 393944
rect 220170 393932 220176 393944
rect 220228 393932 220234 393984
rect 225598 393932 225604 393984
rect 225656 393972 225662 393984
rect 226242 393972 226248 393984
rect 225656 393944 226248 393972
rect 225656 393932 225662 393944
rect 226242 393932 226248 393944
rect 226300 393932 226306 393984
rect 226610 393932 226616 393984
rect 226668 393972 226674 393984
rect 226978 393972 226984 393984
rect 226668 393944 226984 393972
rect 226668 393932 226674 393944
rect 226978 393932 226984 393944
rect 227036 393932 227042 393984
rect 227806 393932 227812 393984
rect 227864 393972 227870 393984
rect 227990 393972 227996 393984
rect 227864 393944 227996 393972
rect 227864 393932 227870 393944
rect 227990 393932 227996 393944
rect 228048 393932 228054 393984
rect 228082 393932 228088 393984
rect 228140 393972 228146 393984
rect 228818 393972 228824 393984
rect 228140 393944 228824 393972
rect 228140 393932 228146 393944
rect 228818 393932 228824 393944
rect 228876 393932 228882 393984
rect 229278 393932 229284 393984
rect 229336 393972 229342 393984
rect 230106 393972 230112 393984
rect 229336 393944 230112 393972
rect 229336 393932 229342 393944
rect 230106 393932 230112 393944
rect 230164 393932 230170 393984
rect 230750 393932 230756 393984
rect 230808 393972 230814 393984
rect 230934 393972 230940 393984
rect 230808 393944 230940 393972
rect 230808 393932 230814 393944
rect 230934 393932 230940 393944
rect 230992 393932 230998 393984
rect 231854 393932 231860 393984
rect 231912 393972 231918 393984
rect 232406 393972 232412 393984
rect 231912 393944 232412 393972
rect 231912 393932 231918 393944
rect 232406 393932 232412 393944
rect 232464 393932 232470 393984
rect 233510 393932 233516 393984
rect 233568 393972 233574 393984
rect 233786 393972 233792 393984
rect 233568 393944 233792 393972
rect 233568 393932 233574 393944
rect 233786 393932 233792 393944
rect 233844 393932 233850 393984
rect 236086 393932 236092 393984
rect 236144 393972 236150 393984
rect 236638 393972 236644 393984
rect 236144 393944 236644 393972
rect 236144 393932 236150 393944
rect 236638 393932 236644 393944
rect 236696 393932 236702 393984
rect 237466 393932 237472 393984
rect 237524 393972 237530 393984
rect 238018 393972 238024 393984
rect 237524 393944 238024 393972
rect 237524 393932 237530 393944
rect 238018 393932 238024 393944
rect 238076 393932 238082 393984
rect 238754 393932 238760 393984
rect 238812 393972 238818 393984
rect 239398 393972 239404 393984
rect 238812 393944 239404 393972
rect 238812 393932 238818 393944
rect 239398 393932 239404 393944
rect 239456 393932 239462 393984
rect 240410 393932 240416 393984
rect 240468 393972 240474 393984
rect 240870 393972 240876 393984
rect 240468 393944 240876 393972
rect 240468 393932 240474 393944
rect 240870 393932 240876 393944
rect 240928 393932 240934 393984
rect 241790 393932 241796 393984
rect 241848 393972 241854 393984
rect 242342 393972 242348 393984
rect 241848 393944 242348 393972
rect 241848 393932 241854 393944
rect 242342 393932 242348 393944
rect 242400 393932 242406 393984
rect 242986 393932 242992 393984
rect 243044 393972 243050 393984
rect 243262 393972 243268 393984
rect 243044 393944 243268 393972
rect 243044 393932 243050 393944
rect 243262 393932 243268 393944
rect 243320 393932 243326 393984
rect 243906 393932 243912 393984
rect 243964 393972 243970 393984
rect 379514 393972 379520 393984
rect 243964 393944 379520 393972
rect 243964 393932 243970 393944
rect 379514 393932 379520 393944
rect 379572 393932 379578 393984
rect 225138 393864 225144 393916
rect 225196 393904 225202 393916
rect 225690 393904 225696 393916
rect 225196 393876 225696 393904
rect 225196 393864 225202 393876
rect 225690 393864 225696 393876
rect 225748 393864 225754 393916
rect 229370 393864 229376 393916
rect 229428 393904 229434 393916
rect 234154 393904 234160 393916
rect 229428 393876 234160 393904
rect 229428 393864 229434 393876
rect 234154 393864 234160 393876
rect 234212 393864 234218 393916
rect 235258 393864 235264 393916
rect 235316 393864 235322 393916
rect 240226 393864 240232 393916
rect 240284 393904 240290 393916
rect 240778 393904 240784 393916
rect 240284 393876 240784 393904
rect 240284 393864 240290 393876
rect 240778 393864 240784 393876
rect 240836 393864 240842 393916
rect 245654 393864 245660 393916
rect 245712 393904 245718 393916
rect 246298 393904 246304 393916
rect 245712 393876 246304 393904
rect 245712 393864 245718 393876
rect 246298 393864 246304 393876
rect 246356 393864 246362 393916
rect 247218 393864 247224 393916
rect 247276 393904 247282 393916
rect 247276 393876 247448 393904
rect 247276 393864 247282 393876
rect 225506 393796 225512 393848
rect 225564 393836 225570 393848
rect 226150 393836 226156 393848
rect 225564 393808 226156 393836
rect 225564 393796 225570 393808
rect 226150 393796 226156 393808
rect 226208 393796 226214 393848
rect 229278 393796 229284 393848
rect 229336 393836 229342 393848
rect 229554 393836 229560 393848
rect 229336 393808 229560 393836
rect 229336 393796 229342 393808
rect 229554 393796 229560 393808
rect 229612 393796 229618 393848
rect 230566 393796 230572 393848
rect 230624 393836 230630 393848
rect 231118 393836 231124 393848
rect 230624 393808 231124 393836
rect 230624 393796 230630 393808
rect 231118 393796 231124 393808
rect 231176 393796 231182 393848
rect 231854 393796 231860 393848
rect 231912 393836 231918 393848
rect 232682 393836 232688 393848
rect 231912 393808 232688 393836
rect 231912 393796 231918 393808
rect 232682 393796 232688 393808
rect 232740 393796 232746 393848
rect 233234 393796 233240 393848
rect 233292 393836 233298 393848
rect 233510 393836 233516 393848
rect 233292 393808 233516 393836
rect 233292 393796 233298 393808
rect 233510 393796 233516 393808
rect 233568 393796 233574 393848
rect 225230 393728 225236 393780
rect 225288 393768 225294 393780
rect 226058 393768 226064 393780
rect 225288 393740 226064 393768
rect 225288 393728 225294 393740
rect 226058 393728 226064 393740
rect 226116 393728 226122 393780
rect 230658 393728 230664 393780
rect 230716 393768 230722 393780
rect 231394 393768 231400 393780
rect 230716 393740 231400 393768
rect 230716 393728 230722 393740
rect 231394 393728 231400 393740
rect 231452 393728 231458 393780
rect 232038 393728 232044 393780
rect 232096 393768 232102 393780
rect 232774 393768 232780 393780
rect 232096 393740 232780 393768
rect 232096 393728 232102 393740
rect 232774 393728 232780 393740
rect 232832 393728 232838 393780
rect 235276 393768 235304 393864
rect 238846 393796 238852 393848
rect 238904 393836 238910 393848
rect 239122 393836 239128 393848
rect 238904 393808 239128 393836
rect 238904 393796 238910 393808
rect 239122 393796 239128 393808
rect 239180 393796 239186 393848
rect 240318 393796 240324 393848
rect 240376 393836 240382 393848
rect 241054 393836 241060 393848
rect 240376 393808 241060 393836
rect 240376 393796 240382 393808
rect 241054 393796 241060 393808
rect 241112 393796 241118 393848
rect 241606 393796 241612 393848
rect 241664 393836 241670 393848
rect 242434 393836 242440 393848
rect 241664 393808 242440 393836
rect 241664 393796 241670 393808
rect 242434 393796 242440 393808
rect 242492 393796 242498 393848
rect 243078 393796 243084 393848
rect 243136 393836 243142 393848
rect 243446 393836 243452 393848
rect 243136 393808 243452 393836
rect 243136 393796 243142 393808
rect 243446 393796 243452 393808
rect 243504 393796 243510 393848
rect 245838 393796 245844 393848
rect 245896 393836 245902 393848
rect 246574 393836 246580 393848
rect 245896 393808 246580 393836
rect 245896 393796 245902 393808
rect 246574 393796 246580 393808
rect 246632 393796 246638 393848
rect 234908 393740 235304 393768
rect 234908 393712 234936 393740
rect 243262 393728 243268 393780
rect 243320 393768 243326 393780
rect 243630 393768 243636 393780
rect 243320 393740 243636 393768
rect 243320 393728 243326 393740
rect 243630 393728 243636 393740
rect 243688 393728 243694 393780
rect 245930 393728 245936 393780
rect 245988 393768 245994 393780
rect 246114 393768 246120 393780
rect 245988 393740 246120 393768
rect 245988 393728 245994 393740
rect 246114 393728 246120 393740
rect 246172 393728 246178 393780
rect 247420 393712 247448 393876
rect 248414 393864 248420 393916
rect 248472 393904 248478 393916
rect 248782 393904 248788 393916
rect 248472 393876 248788 393904
rect 248472 393864 248478 393876
rect 248782 393864 248788 393876
rect 248840 393864 248846 393916
rect 249794 393864 249800 393916
rect 249852 393904 249858 393916
rect 250162 393904 250168 393916
rect 249852 393876 250168 393904
rect 249852 393864 249858 393876
rect 250162 393864 250168 393876
rect 250220 393864 250226 393916
rect 250254 393864 250260 393916
rect 250312 393904 250318 393916
rect 250622 393904 250628 393916
rect 250312 393876 250628 393904
rect 250312 393864 250318 393876
rect 250622 393864 250628 393876
rect 250680 393864 250686 393916
rect 251726 393864 251732 393916
rect 251784 393904 251790 393916
rect 251910 393904 251916 393916
rect 251784 393876 251916 393904
rect 251784 393864 251790 393876
rect 251910 393864 251916 393876
rect 251968 393864 251974 393916
rect 254578 393864 254584 393916
rect 254636 393904 254642 393916
rect 254946 393904 254952 393916
rect 254636 393876 254952 393904
rect 254636 393864 254642 393876
rect 254946 393864 254952 393876
rect 255004 393864 255010 393916
rect 251358 393796 251364 393848
rect 251416 393836 251422 393848
rect 251634 393836 251640 393848
rect 251416 393808 251640 393836
rect 251416 393796 251422 393808
rect 251634 393796 251640 393808
rect 251692 393796 251698 393848
rect 252646 393796 252652 393848
rect 252704 393836 252710 393848
rect 252830 393836 252836 393848
rect 252704 393808 252836 393836
rect 252704 393796 252710 393808
rect 252830 393796 252836 393808
rect 252888 393796 252894 393848
rect 253014 393796 253020 393848
rect 253072 393836 253078 393848
rect 253382 393836 253388 393848
rect 253072 393808 253388 393836
rect 253072 393796 253078 393808
rect 253382 393796 253388 393808
rect 253440 393796 253446 393848
rect 254302 393796 254308 393848
rect 254360 393836 254366 393848
rect 254486 393836 254492 393848
rect 254360 393808 254492 393836
rect 254360 393796 254366 393808
rect 254486 393796 254492 393808
rect 254544 393796 254550 393848
rect 255314 393796 255320 393848
rect 255372 393836 255378 393848
rect 255590 393836 255596 393848
rect 255372 393808 255596 393836
rect 255372 393796 255378 393808
rect 255590 393796 255596 393808
rect 255648 393796 255654 393848
rect 248414 393728 248420 393780
rect 248472 393768 248478 393780
rect 249334 393768 249340 393780
rect 248472 393740 249340 393768
rect 248472 393728 248478 393740
rect 249334 393728 249340 393740
rect 249392 393728 249398 393780
rect 251266 393728 251272 393780
rect 251324 393768 251330 393780
rect 252094 393768 252100 393780
rect 251324 393740 252100 393768
rect 251324 393728 251330 393740
rect 252094 393728 252100 393740
rect 252152 393728 252158 393780
rect 254210 393728 254216 393780
rect 254268 393768 254274 393780
rect 254670 393768 254676 393780
rect 254268 393740 254676 393768
rect 254268 393728 254274 393740
rect 254670 393728 254676 393740
rect 254728 393728 254734 393780
rect 226426 393660 226432 393712
rect 226484 393700 226490 393712
rect 227070 393700 227076 393712
rect 226484 393672 227076 393700
rect 226484 393660 226490 393672
rect 227070 393660 227076 393672
rect 227128 393660 227134 393712
rect 227990 393660 227996 393712
rect 228048 393700 228054 393712
rect 228358 393700 228364 393712
rect 228048 393672 228364 393700
rect 228048 393660 228054 393672
rect 228358 393660 228364 393672
rect 228416 393660 228422 393712
rect 230842 393660 230848 393712
rect 230900 393700 230906 393712
rect 231210 393700 231216 393712
rect 230900 393672 231216 393700
rect 230900 393660 230906 393672
rect 231210 393660 231216 393672
rect 231268 393660 231274 393712
rect 234890 393660 234896 393712
rect 234948 393660 234954 393712
rect 235074 393660 235080 393712
rect 235132 393700 235138 393712
rect 235442 393700 235448 393712
rect 235132 393672 235448 393700
rect 235132 393660 235138 393672
rect 235442 393660 235448 393672
rect 235500 393660 235506 393712
rect 243078 393660 243084 393712
rect 243136 393700 243142 393712
rect 243814 393700 243820 393712
rect 243136 393672 243820 393700
rect 243136 393660 243142 393672
rect 243814 393660 243820 393672
rect 243872 393660 243878 393712
rect 244366 393660 244372 393712
rect 244424 393700 244430 393712
rect 245194 393700 245200 393712
rect 244424 393672 245200 393700
rect 244424 393660 244430 393672
rect 245194 393660 245200 393672
rect 245252 393660 245258 393712
rect 247402 393660 247408 393712
rect 247460 393660 247466 393712
rect 248690 393660 248696 393712
rect 248748 393700 248754 393712
rect 249150 393700 249156 393712
rect 248748 393672 249156 393700
rect 248748 393660 248754 393672
rect 249150 393660 249156 393672
rect 249208 393660 249214 393712
rect 252462 393660 252468 393712
rect 252520 393700 252526 393712
rect 253106 393700 253112 393712
rect 252520 393672 253112 393700
rect 252520 393660 252526 393672
rect 253106 393660 253112 393672
rect 253164 393660 253170 393712
rect 254026 393660 254032 393712
rect 254084 393700 254090 393712
rect 254486 393700 254492 393712
rect 254084 393672 254492 393700
rect 254084 393660 254090 393672
rect 254486 393660 254492 393672
rect 254544 393660 254550 393712
rect 226886 393592 226892 393644
rect 226944 393632 226950 393644
rect 227622 393632 227628 393644
rect 226944 393604 227628 393632
rect 226944 393592 226950 393604
rect 227622 393592 227628 393604
rect 227680 393592 227686 393644
rect 227714 393592 227720 393644
rect 227772 393632 227778 393644
rect 228082 393632 228088 393644
rect 227772 393604 228088 393632
rect 227772 393592 227778 393604
rect 228082 393592 228088 393604
rect 228140 393592 228146 393644
rect 246114 393592 246120 393644
rect 246172 393632 246178 393644
rect 246390 393632 246396 393644
rect 246172 393604 246396 393632
rect 246172 393592 246178 393604
rect 246390 393592 246396 393604
rect 246448 393592 246454 393644
rect 227898 393524 227904 393576
rect 227956 393564 227962 393576
rect 228450 393564 228456 393576
rect 227956 393536 228456 393564
rect 227956 393524 227962 393536
rect 228450 393524 228456 393536
rect 228508 393524 228514 393576
rect 230382 393524 230388 393576
rect 230440 393564 230446 393576
rect 231210 393564 231216 393576
rect 230440 393536 231216 393564
rect 230440 393524 230446 393536
rect 231210 393524 231216 393536
rect 231268 393524 231274 393576
rect 239122 393524 239128 393576
rect 239180 393564 239186 393576
rect 239582 393564 239588 393576
rect 239180 393536 239588 393564
rect 239180 393524 239186 393536
rect 239582 393524 239588 393536
rect 239640 393524 239646 393576
rect 254026 393524 254032 393576
rect 254084 393564 254090 393576
rect 254854 393564 254860 393576
rect 254084 393536 254860 393564
rect 254084 393524 254090 393536
rect 254854 393524 254860 393536
rect 254912 393524 254918 393576
rect 236270 393456 236276 393508
rect 236328 393496 236334 393508
rect 236454 393496 236460 393508
rect 236328 393468 236460 393496
rect 236328 393456 236334 393468
rect 236454 393456 236460 393468
rect 236512 393456 236518 393508
rect 239030 393456 239036 393508
rect 239088 393496 239094 393508
rect 239490 393496 239496 393508
rect 239088 393468 239496 393496
rect 239088 393456 239094 393468
rect 239490 393456 239496 393468
rect 239548 393456 239554 393508
rect 231486 392844 231492 392896
rect 231544 392884 231550 392896
rect 257614 392884 257620 392896
rect 231544 392856 257620 392884
rect 231544 392844 231550 392856
rect 257614 392844 257620 392856
rect 257672 392844 257678 392896
rect 232866 392776 232872 392828
rect 232924 392816 232930 392828
rect 277394 392816 277400 392828
rect 232924 392788 277400 392816
rect 232924 392776 232930 392788
rect 277394 392776 277400 392788
rect 277452 392776 277458 392828
rect 238386 392708 238392 392760
rect 238444 392748 238450 392760
rect 349154 392748 349160 392760
rect 238444 392720 349160 392748
rect 238444 392708 238450 392720
rect 349154 392708 349160 392720
rect 349212 392708 349218 392760
rect 164234 392640 164240 392692
rect 164292 392680 164298 392692
rect 215938 392680 215944 392692
rect 164292 392652 215944 392680
rect 164292 392640 164298 392652
rect 215938 392640 215944 392652
rect 215996 392640 216002 392692
rect 245010 392640 245016 392692
rect 245068 392680 245074 392692
rect 445754 392680 445760 392692
rect 245068 392652 445760 392680
rect 245068 392640 245074 392652
rect 445754 392640 445760 392652
rect 445812 392640 445818 392692
rect 34514 392572 34520 392624
rect 34572 392612 34578 392624
rect 213362 392612 213368 392624
rect 34572 392584 213368 392612
rect 34572 392572 34578 392584
rect 213362 392572 213368 392584
rect 213420 392572 213426 392624
rect 248046 392572 248052 392624
rect 248104 392612 248110 392624
rect 480254 392612 480260 392624
rect 248104 392584 480260 392612
rect 248104 392572 248110 392584
rect 480254 392572 480260 392584
rect 480312 392572 480318 392624
rect 249978 392300 249984 392352
rect 250036 392340 250042 392352
rect 250530 392340 250536 392352
rect 250036 392312 250536 392340
rect 250036 392300 250042 392312
rect 250530 392300 250536 392312
rect 250588 392300 250594 392352
rect 251174 392300 251180 392352
rect 251232 392340 251238 392352
rect 251818 392340 251824 392352
rect 251232 392312 251824 392340
rect 251232 392300 251238 392312
rect 251818 392300 251824 392312
rect 251876 392300 251882 392352
rect 229186 392164 229192 392216
rect 229244 392204 229250 392216
rect 229462 392204 229468 392216
rect 229244 392176 229468 392204
rect 229244 392164 229250 392176
rect 229462 392164 229468 392176
rect 229520 392164 229526 392216
rect 233418 392164 233424 392216
rect 233476 392204 233482 392216
rect 233694 392204 233700 392216
rect 233476 392176 233700 392204
rect 233476 392164 233482 392176
rect 233694 392164 233700 392176
rect 233752 392164 233758 392216
rect 237558 392164 237564 392216
rect 237616 392204 237622 392216
rect 237742 392204 237748 392216
rect 237616 392176 237748 392204
rect 237616 392164 237622 392176
rect 237742 392164 237748 392176
rect 237800 392164 237806 392216
rect 233326 392096 233332 392148
rect 233384 392136 233390 392148
rect 233878 392136 233884 392148
rect 233384 392108 233884 392136
rect 233384 392096 233390 392108
rect 233878 392096 233884 392108
rect 233936 392096 233942 392148
rect 229094 392028 229100 392080
rect 229152 392068 229158 392080
rect 229738 392068 229744 392080
rect 229152 392040 229744 392068
rect 229152 392028 229158 392040
rect 229738 392028 229744 392040
rect 229796 392028 229802 392080
rect 237558 392028 237564 392080
rect 237616 392068 237622 392080
rect 238294 392068 238300 392080
rect 237616 392040 238300 392068
rect 237616 392028 237622 392040
rect 238294 392028 238300 392040
rect 238352 392028 238358 392080
rect 229278 391892 229284 391944
rect 229336 391932 229342 391944
rect 230014 391932 230020 391944
rect 229336 391904 230020 391932
rect 229336 391892 229342 391904
rect 230014 391892 230020 391904
rect 230072 391892 230078 391944
rect 228726 391824 228732 391876
rect 228784 391864 228790 391876
rect 233510 391864 233516 391876
rect 228784 391836 233516 391864
rect 228784 391824 228790 391836
rect 233510 391824 233516 391836
rect 233568 391824 233574 391876
rect 225414 391688 225420 391740
rect 225472 391728 225478 391740
rect 225966 391728 225972 391740
rect 225472 391700 225972 391728
rect 225472 391688 225478 391700
rect 225966 391688 225972 391700
rect 226024 391688 226030 391740
rect 240042 391484 240048 391536
rect 240100 391524 240106 391536
rect 313274 391524 313280 391536
rect 240100 391496 313280 391524
rect 240100 391484 240106 391496
rect 313274 391484 313280 391496
rect 313332 391484 313338 391536
rect 240962 391416 240968 391468
rect 241020 391456 241026 391468
rect 385034 391456 385040 391468
rect 241020 391428 385040 391456
rect 241020 391416 241026 391428
rect 385034 391416 385040 391428
rect 385092 391416 385098 391468
rect 243722 391348 243728 391400
rect 243780 391388 243786 391400
rect 419534 391388 419540 391400
rect 243780 391360 419540 391388
rect 243780 391348 243786 391360
rect 419534 391348 419540 391360
rect 419592 391348 419598 391400
rect 236362 391280 236368 391332
rect 236420 391320 236426 391332
rect 236420 391292 236500 391320
rect 236420 391280 236426 391292
rect 184934 391212 184940 391264
rect 184992 391252 184998 391264
rect 224310 391252 224316 391264
rect 184992 391224 224316 391252
rect 184992 391212 184998 391224
rect 224310 391212 224316 391224
rect 224368 391212 224374 391264
rect 236472 391128 236500 391292
rect 245378 391280 245384 391332
rect 245436 391320 245442 391332
rect 437474 391320 437480 391332
rect 245436 391292 437480 391320
rect 245436 391280 245442 391292
rect 437474 391280 437480 391292
rect 437532 391280 437538 391332
rect 249242 391212 249248 391264
rect 249300 391252 249306 391264
rect 492674 391252 492680 391264
rect 249300 391224 492680 391252
rect 249300 391212 249306 391224
rect 492674 391212 492680 391224
rect 492732 391212 492738 391264
rect 236454 391076 236460 391128
rect 236512 391076 236518 391128
rect 252830 391008 252836 391060
rect 252888 391048 252894 391060
rect 253290 391048 253296 391060
rect 252888 391020 253296 391048
rect 252888 391008 252894 391020
rect 253290 391008 253296 391020
rect 253348 391008 253354 391060
rect 247310 390396 247316 390448
rect 247368 390436 247374 390448
rect 247770 390436 247776 390448
rect 247368 390408 247776 390436
rect 247368 390396 247374 390408
rect 247770 390396 247776 390408
rect 247828 390396 247834 390448
rect 247586 390328 247592 390380
rect 247644 390368 247650 390380
rect 247644 390340 247816 390368
rect 247644 390328 247650 390340
rect 247788 390176 247816 390340
rect 247770 390124 247776 390176
rect 247828 390124 247834 390176
rect 234062 389784 234068 389836
rect 234120 389824 234126 389836
rect 300854 389824 300860 389836
rect 234120 389796 300860 389824
rect 234120 389784 234126 389796
rect 300854 389784 300860 389796
rect 300912 389784 300918 389836
rect 233510 389376 233516 389428
rect 233568 389416 233574 389428
rect 233970 389416 233976 389428
rect 233568 389388 233976 389416
rect 233568 389376 233574 389388
rect 233970 389376 233976 389388
rect 234028 389376 234034 389428
rect 233418 389240 233424 389292
rect 233476 389240 233482 389292
rect 233436 389212 233464 389240
rect 233786 389212 233792 389224
rect 233436 389184 233792 389212
rect 233786 389172 233792 389184
rect 233844 389172 233850 389224
rect 233878 389172 233884 389224
rect 233936 389212 233942 389224
rect 234154 389212 234160 389224
rect 233936 389184 234160 389212
rect 233936 389172 233942 389184
rect 234154 389172 234160 389184
rect 234212 389172 234218 389224
rect 227162 386520 227168 386572
rect 227220 386560 227226 386572
rect 227530 386560 227536 386572
rect 227220 386532 227536 386560
rect 227220 386520 227226 386532
rect 227530 386520 227536 386532
rect 227588 386520 227594 386572
rect 299106 379448 299112 379500
rect 299164 379488 299170 379500
rect 580166 379488 580172 379500
rect 299164 379460 580172 379488
rect 299164 379448 299170 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3050 372512 3056 372564
rect 3108 372552 3114 372564
rect 106918 372552 106924 372564
rect 3108 372524 106924 372552
rect 3108 372512 3114 372524
rect 106918 372512 106924 372524
rect 106976 372512 106982 372564
rect 296622 365644 296628 365696
rect 296680 365684 296686 365696
rect 580166 365684 580172 365696
rect 296680 365656 580172 365684
rect 296680 365644 296686 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3510 358708 3516 358760
rect 3568 358748 3574 358760
rect 184198 358748 184204 358760
rect 3568 358720 184204 358748
rect 3568 358708 3574 358720
rect 184198 358708 184204 358720
rect 184256 358708 184262 358760
rect 23474 358028 23480 358080
rect 23532 358068 23538 358080
rect 208210 358068 208216 358080
rect 23532 358040 208216 358068
rect 23532 358028 23538 358040
rect 208210 358028 208216 358040
rect 208268 358028 208274 358080
rect 237926 356668 237932 356720
rect 237984 356708 237990 356720
rect 350534 356708 350540 356720
rect 237984 356680 350540 356708
rect 237984 356668 237990 356680
rect 350534 356668 350540 356680
rect 350592 356668 350598 356720
rect 235258 355648 235264 355700
rect 235316 355688 235322 355700
rect 316034 355688 316040 355700
rect 235316 355660 316040 355688
rect 235316 355648 235322 355660
rect 316034 355648 316040 355660
rect 316092 355648 316098 355700
rect 235442 355580 235448 355632
rect 235500 355620 235506 355632
rect 324406 355620 324412 355632
rect 235500 355592 324412 355620
rect 235500 355580 235506 355592
rect 324406 355580 324412 355592
rect 324464 355580 324470 355632
rect 113174 355512 113180 355564
rect 113232 355552 113238 355564
rect 218698 355552 218704 355564
rect 113232 355524 218704 355552
rect 113232 355512 113238 355524
rect 218698 355512 218704 355524
rect 218756 355512 218762 355564
rect 242434 355512 242440 355564
rect 242492 355552 242498 355564
rect 357434 355552 357440 355564
rect 242492 355524 357440 355552
rect 242492 355512 242498 355524
rect 357434 355512 357440 355524
rect 357492 355512 357498 355564
rect 88334 355444 88340 355496
rect 88392 355484 88398 355496
rect 213270 355484 213276 355496
rect 88392 355456 213276 355484
rect 88392 355444 88398 355456
rect 213270 355444 213276 355456
rect 213328 355444 213334 355496
rect 239214 355444 239220 355496
rect 239272 355484 239278 355496
rect 367094 355484 367100 355496
rect 239272 355456 367100 355484
rect 239272 355444 239278 355456
rect 367094 355444 367100 355456
rect 367152 355444 367158 355496
rect 73154 355376 73160 355428
rect 73212 355416 73218 355428
rect 215846 355416 215852 355428
rect 73212 355388 215852 355416
rect 73212 355376 73218 355388
rect 215846 355376 215852 355388
rect 215904 355376 215910 355428
rect 239306 355376 239312 355428
rect 239364 355416 239370 355428
rect 371234 355416 371240 355428
rect 239364 355388 371240 355416
rect 239364 355376 239370 355388
rect 371234 355376 371240 355388
rect 371292 355376 371298 355428
rect 45554 355308 45560 355360
rect 45612 355348 45618 355360
rect 204990 355348 204996 355360
rect 45612 355320 204996 355348
rect 45612 355308 45618 355320
rect 204990 355308 204996 355320
rect 205048 355308 205054 355360
rect 246666 355308 246672 355360
rect 246724 355348 246730 355360
rect 393314 355348 393320 355360
rect 246724 355320 393320 355348
rect 246724 355308 246730 355320
rect 393314 355308 393320 355320
rect 393372 355308 393378 355360
rect 78674 354356 78680 354408
rect 78732 354396 78738 354408
rect 215754 354396 215760 354408
rect 78732 354368 215760 354396
rect 78732 354356 78738 354368
rect 215754 354356 215760 354368
rect 215812 354356 215818 354408
rect 56594 354288 56600 354340
rect 56652 354328 56658 354340
rect 211890 354328 211896 354340
rect 56652 354300 211896 354328
rect 56652 354288 56658 354300
rect 211890 354288 211896 354300
rect 211948 354288 211954 354340
rect 231302 354288 231308 354340
rect 231360 354328 231366 354340
rect 269114 354328 269120 354340
rect 231360 354300 269120 354328
rect 231360 354288 231366 354300
rect 269114 354288 269120 354300
rect 269172 354288 269178 354340
rect 42794 354220 42800 354272
rect 42852 354260 42858 354272
rect 212994 354260 213000 354272
rect 42852 354232 213000 354260
rect 42852 354220 42858 354232
rect 212994 354220 213000 354232
rect 213052 354220 213058 354272
rect 232590 354220 232596 354272
rect 232648 354260 232654 354272
rect 284294 354260 284300 354272
rect 232648 354232 284300 354260
rect 232648 354220 232654 354232
rect 284294 354220 284300 354232
rect 284352 354220 284358 354272
rect 41414 354152 41420 354204
rect 41472 354192 41478 354204
rect 212902 354192 212908 354204
rect 41472 354164 212908 354192
rect 41472 354152 41478 354164
rect 212902 354152 212908 354164
rect 212960 354152 212966 354204
rect 238018 354152 238024 354204
rect 238076 354192 238082 354204
rect 357526 354192 357532 354204
rect 238076 354164 357532 354192
rect 238076 354152 238082 354164
rect 357526 354152 357532 354164
rect 357584 354152 357590 354204
rect 19334 354084 19340 354136
rect 19392 354124 19398 354136
rect 211614 354124 211620 354136
rect 19392 354096 211620 354124
rect 19392 354084 19398 354096
rect 211614 354084 211620 354096
rect 211672 354084 211678 354136
rect 240778 354084 240784 354136
rect 240836 354124 240842 354136
rect 397454 354124 397460 354136
rect 240836 354096 397460 354124
rect 240836 354084 240842 354096
rect 397454 354084 397460 354096
rect 397512 354084 397518 354136
rect 19426 354016 19432 354068
rect 19484 354056 19490 354068
rect 211706 354056 211712 354068
rect 19484 354028 211712 354056
rect 19484 354016 19490 354028
rect 211706 354016 211712 354028
rect 211764 354016 211770 354068
rect 229738 354016 229744 354068
rect 229796 354056 229802 354068
rect 242066 354056 242072 354068
rect 229796 354028 242072 354056
rect 229796 354016 229802 354028
rect 242066 354016 242072 354028
rect 242124 354016 242130 354068
rect 251910 354016 251916 354068
rect 251968 354056 251974 354068
rect 531314 354056 531320 354068
rect 251968 354028 531320 354056
rect 251968 354016 251974 354028
rect 531314 354016 531320 354028
rect 531372 354016 531378 354068
rect 13814 353948 13820 354000
rect 13872 353988 13878 354000
rect 210694 353988 210700 354000
rect 13872 353960 210700 353988
rect 13872 353948 13878 353960
rect 210694 353948 210700 353960
rect 210752 353948 210758 354000
rect 229830 353948 229836 354000
rect 229888 353988 229894 354000
rect 251634 353988 251640 354000
rect 229888 353960 251640 353988
rect 229888 353948 229894 353960
rect 251634 353948 251640 353960
rect 251692 353948 251698 354000
rect 254670 353948 254676 354000
rect 254728 353988 254734 354000
rect 560294 353988 560300 354000
rect 254728 353960 560300 353988
rect 254728 353948 254734 353960
rect 560294 353948 560300 353960
rect 560352 353948 560358 354000
rect 231210 352792 231216 352844
rect 231268 352832 231274 352844
rect 259546 352832 259552 352844
rect 231268 352804 259552 352832
rect 231268 352792 231274 352804
rect 259546 352792 259552 352804
rect 259604 352792 259610 352844
rect 157334 352724 157340 352776
rect 157392 352764 157398 352776
rect 222746 352764 222752 352776
rect 157392 352736 222752 352764
rect 157392 352724 157398 352736
rect 222746 352724 222752 352736
rect 222804 352724 222810 352776
rect 231026 352724 231032 352776
rect 231084 352764 231090 352776
rect 266354 352764 266360 352776
rect 231084 352736 266360 352764
rect 231084 352724 231090 352736
rect 266354 352724 266360 352736
rect 266412 352724 266418 352776
rect 104894 352656 104900 352708
rect 104952 352696 104958 352708
rect 218606 352696 218612 352708
rect 104952 352668 218612 352696
rect 104952 352656 104958 352668
rect 218606 352656 218612 352668
rect 218664 352656 218670 352708
rect 257706 352656 257712 352708
rect 257764 352696 257770 352708
rect 436094 352696 436100 352708
rect 257764 352668 436100 352696
rect 257764 352656 257770 352668
rect 436094 352656 436100 352668
rect 436152 352656 436158 352708
rect 52454 352588 52460 352640
rect 52512 352628 52518 352640
rect 214650 352628 214656 352640
rect 52512 352600 214656 352628
rect 52512 352588 52518 352600
rect 214650 352588 214656 352600
rect 214708 352588 214714 352640
rect 250530 352588 250536 352640
rect 250588 352628 250594 352640
rect 511994 352628 512000 352640
rect 250588 352600 512000 352628
rect 250588 352588 250594 352600
rect 511994 352588 512000 352600
rect 512052 352588 512058 352640
rect 3510 352520 3516 352572
rect 3568 352560 3574 352572
rect 201954 352560 201960 352572
rect 3568 352532 201960 352560
rect 3568 352520 3574 352532
rect 201954 352520 201960 352532
rect 202012 352520 202018 352572
rect 213270 352520 213276 352572
rect 213328 352560 213334 352572
rect 227070 352560 227076 352572
rect 213328 352532 227076 352560
rect 213328 352520 213334 352532
rect 227070 352520 227076 352532
rect 227128 352520 227134 352572
rect 228358 352520 228364 352572
rect 228416 352560 228422 352572
rect 235258 352560 235264 352572
rect 228416 352532 235264 352560
rect 228416 352520 228422 352532
rect 235258 352520 235264 352532
rect 235316 352520 235322 352572
rect 251818 352520 251824 352572
rect 251876 352560 251882 352572
rect 524414 352560 524420 352572
rect 251876 352532 524420 352560
rect 251876 352520 251882 352532
rect 524414 352520 524420 352532
rect 524472 352520 524478 352572
rect 204254 351364 204260 351416
rect 204312 351404 204318 351416
rect 225598 351404 225604 351416
rect 204312 351376 225604 351404
rect 204312 351364 204318 351376
rect 225598 351364 225604 351376
rect 225656 351364 225662 351416
rect 182174 351296 182180 351348
rect 182232 351336 182238 351348
rect 224126 351336 224132 351348
rect 182232 351308 224132 351336
rect 182232 351296 182238 351308
rect 224126 351296 224132 351308
rect 224184 351296 224190 351348
rect 151906 351228 151912 351280
rect 151964 351268 151970 351280
rect 221366 351268 221372 351280
rect 151964 351240 221372 351268
rect 151964 351228 151970 351240
rect 221366 351228 221372 351240
rect 221424 351228 221430 351280
rect 236546 351228 236552 351280
rect 236604 351268 236610 351280
rect 342254 351268 342260 351280
rect 236604 351240 342260 351268
rect 236604 351228 236610 351240
rect 342254 351228 342260 351240
rect 342312 351228 342318 351280
rect 4154 351160 4160 351212
rect 4212 351200 4218 351212
rect 209314 351200 209320 351212
rect 4212 351172 209320 351200
rect 4212 351160 4218 351172
rect 209314 351160 209320 351172
rect 209372 351160 209378 351212
rect 253290 351160 253296 351212
rect 253348 351200 253354 351212
rect 554774 351200 554780 351212
rect 253348 351172 554780 351200
rect 253348 351160 253354 351172
rect 554774 351160 554780 351172
rect 554832 351160 554838 351212
rect 222746 350548 222752 350600
rect 222804 350588 222810 350600
rect 226886 350588 226892 350600
rect 222804 350560 226892 350588
rect 222804 350548 222810 350560
rect 226886 350548 226892 350560
rect 226944 350548 226950 350600
rect 254578 347012 254584 347064
rect 254636 347052 254642 347064
rect 572714 347052 572720 347064
rect 254636 347024 572720 347052
rect 254636 347012 254642 347024
rect 572714 347012 572720 347024
rect 572772 347012 572778 347064
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 202046 346372 202052 346384
rect 3200 346344 202052 346372
rect 3200 346332 3206 346344
rect 202046 346332 202052 346344
rect 202104 346332 202110 346384
rect 260190 335996 260196 336048
rect 260248 336036 260254 336048
rect 460934 336036 460940 336048
rect 260248 336008 460940 336036
rect 260248 335996 260254 336008
rect 460934 335996 460940 336008
rect 460992 335996 460998 336048
rect 299014 325592 299020 325644
rect 299072 325632 299078 325644
rect 579890 325632 579896 325644
rect 299072 325604 579896 325632
rect 299072 325592 299078 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 2774 320084 2780 320136
rect 2832 320124 2838 320136
rect 6270 320124 6276 320136
rect 2832 320096 6276 320124
rect 2832 320084 2838 320096
rect 6270 320084 6276 320096
rect 6328 320084 6334 320136
rect 296530 313216 296536 313268
rect 296588 313256 296594 313268
rect 580166 313256 580172 313268
rect 296588 313228 580172 313256
rect 296588 313216 296594 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 14458 306320 14464 306332
rect 3384 306292 14464 306320
rect 3384 306280 3390 306292
rect 14458 306280 14464 306292
rect 14516 306280 14522 306332
rect 258810 302880 258816 302932
rect 258868 302920 258874 302932
rect 449894 302920 449900 302932
rect 258868 302892 449900 302920
rect 258868 302880 258874 302892
rect 449894 302880 449900 302892
rect 449952 302880 449958 302932
rect 3234 293904 3240 293956
rect 3292 293944 3298 293956
rect 202782 293944 202788 293956
rect 3292 293916 202788 293944
rect 3292 293904 3298 293916
rect 202782 293904 202788 293916
rect 202840 293904 202846 293956
rect 298922 273164 298928 273216
rect 298980 273204 298986 273216
rect 579890 273204 579896 273216
rect 298980 273176 579896 273204
rect 298980 273164 298986 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 186958 267696 186964 267708
rect 3292 267668 186964 267696
rect 3292 267656 3298 267668
rect 186958 267656 186964 267668
rect 187016 267656 187022 267708
rect 296438 259360 296444 259412
rect 296496 259400 296502 259412
rect 579798 259400 579804 259412
rect 296496 259372 579804 259400
rect 296496 259360 296502 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3142 254736 3148 254788
rect 3200 254776 3206 254788
rect 6178 254776 6184 254788
rect 3200 254748 6184 254776
rect 3200 254736 3206 254748
rect 6178 254736 6184 254748
rect 6236 254736 6242 254788
rect 298830 245556 298836 245608
rect 298888 245596 298894 245608
rect 580166 245596 580172 245608
rect 298888 245568 580172 245596
rect 298888 245556 298894 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3326 241408 3332 241460
rect 3384 241448 3390 241460
rect 191098 241448 191104 241460
rect 3384 241420 191104 241448
rect 3384 241408 3390 241420
rect 191098 241408 191104 241420
rect 191156 241408 191162 241460
rect 265802 233180 265808 233232
rect 265860 233220 265866 233232
rect 580166 233220 580172 233232
rect 265860 233192 580172 233220
rect 265860 233180 265866 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 246298 228352 246304 228404
rect 246356 228392 246362 228404
rect 386414 228392 386420 228404
rect 246356 228364 386420 228392
rect 246356 228352 246362 228364
rect 386414 228352 386420 228364
rect 386472 228352 386478 228404
rect 296346 219376 296352 219428
rect 296404 219416 296410 219428
rect 579890 219416 579896 219428
rect 296404 219388 579896 219416
rect 296404 219376 296410 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 3142 215228 3148 215280
rect 3200 215268 3206 215280
rect 203610 215268 203616 215280
rect 3200 215240 203616 215268
rect 3200 215228 3206 215240
rect 203610 215228 203616 215240
rect 203668 215228 203674 215280
rect 264330 206932 264336 206984
rect 264388 206972 264394 206984
rect 580166 206972 580172 206984
rect 264388 206944 580172 206972
rect 264388 206932 264394 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 202598 202824 202604 202836
rect 3384 202796 202604 202824
rect 3384 202784 3390 202796
rect 202598 202784 202604 202796
rect 202656 202784 202662 202836
rect 298738 193128 298744 193180
rect 298796 193168 298802 193180
rect 580166 193168 580172 193180
rect 298796 193140 580172 193168
rect 298796 193128 298802 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 262858 182792 262864 182844
rect 262916 182832 262922 182844
rect 467834 182832 467840 182844
rect 262916 182804 467840 182832
rect 262916 182792 262922 182804
rect 467834 182792 467840 182804
rect 467892 182792 467898 182844
rect 296254 179324 296260 179376
rect 296312 179364 296318 179376
rect 579982 179364 579988 179376
rect 296312 179336 579988 179364
rect 296312 179324 296318 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 233786 177692 233792 177744
rect 233844 177732 233850 177744
rect 293954 177732 293960 177744
rect 233844 177704 293960 177732
rect 233844 177692 233850 177704
rect 293954 177692 293960 177704
rect 294012 177692 294018 177744
rect 233970 177624 233976 177676
rect 234028 177664 234034 177676
rect 298094 177664 298100 177676
rect 234028 177636 298100 177664
rect 234028 177624 234034 177636
rect 298094 177624 298100 177636
rect 298152 177624 298158 177676
rect 203058 177556 203064 177608
rect 203116 177596 203122 177608
rect 225506 177596 225512 177608
rect 203116 177568 225512 177596
rect 203116 177556 203122 177568
rect 225506 177556 225512 177568
rect 225564 177556 225570 177608
rect 240686 177556 240692 177608
rect 240744 177596 240750 177608
rect 382274 177596 382280 177608
rect 240744 177568 382280 177596
rect 240744 177556 240750 177568
rect 382274 177556 382280 177568
rect 382332 177556 382338 177608
rect 201494 177488 201500 177540
rect 201552 177528 201558 177540
rect 225414 177528 225420 177540
rect 201552 177500 225420 177528
rect 201552 177488 201558 177500
rect 225414 177488 225420 177500
rect 225472 177488 225478 177540
rect 240594 177488 240600 177540
rect 240652 177528 240658 177540
rect 390554 177528 390560 177540
rect 240652 177500 390560 177528
rect 240652 177488 240658 177500
rect 390554 177488 390560 177500
rect 390612 177488 390618 177540
rect 133874 177420 133880 177472
rect 133932 177460 133938 177472
rect 219986 177460 219992 177472
rect 133932 177432 219992 177460
rect 133932 177420 133938 177432
rect 219986 177420 219992 177432
rect 220044 177420 220050 177472
rect 247678 177420 247684 177472
rect 247736 177460 247742 177472
rect 478874 177460 478880 177472
rect 247736 177432 478880 177460
rect 247736 177420 247742 177432
rect 478874 177420 478880 177432
rect 478932 177420 478938 177472
rect 126974 177352 126980 177404
rect 127032 177392 127038 177404
rect 219894 177392 219900 177404
rect 127032 177364 219900 177392
rect 127032 177352 127038 177364
rect 219894 177352 219900 177364
rect 219952 177352 219958 177404
rect 250438 177352 250444 177404
rect 250496 177392 250502 177404
rect 518894 177392 518900 177404
rect 250496 177364 518900 177392
rect 250496 177352 250502 177364
rect 518894 177352 518900 177364
rect 518952 177352 518958 177404
rect 77386 177284 77392 177336
rect 77444 177324 77450 177336
rect 210602 177324 210608 177336
rect 77444 177296 210608 177324
rect 77444 177284 77450 177296
rect 210602 177284 210608 177296
rect 210660 177284 210666 177336
rect 215754 177284 215760 177336
rect 215812 177324 215818 177336
rect 226794 177324 226800 177336
rect 215812 177296 226800 177324
rect 215812 177284 215818 177296
rect 226794 177284 226800 177296
rect 226852 177284 226858 177336
rect 251726 177284 251732 177336
rect 251784 177324 251790 177336
rect 532694 177324 532700 177336
rect 251784 177296 532700 177324
rect 251784 177284 251790 177296
rect 532694 177284 532700 177296
rect 532752 177284 532758 177336
rect 38654 175924 38660 175976
rect 38712 175964 38718 175976
rect 206462 175964 206468 175976
rect 38712 175936 206468 175964
rect 38712 175924 38718 175936
rect 206462 175924 206468 175936
rect 206520 175924 206526 175976
rect 102134 171776 102140 171828
rect 102192 171816 102198 171828
rect 209222 171816 209228 171828
rect 102192 171788 209228 171816
rect 102192 171776 102198 171788
rect 209222 171776 209228 171788
rect 209280 171776 209286 171828
rect 272518 166948 272524 167000
rect 272576 166988 272582 167000
rect 580166 166988 580172 167000
rect 272576 166960 580172 166988
rect 272576 166948 272582 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 199378 164200 199384 164212
rect 3384 164172 199384 164200
rect 3384 164160 3390 164172
rect 199378 164160 199384 164172
rect 199436 164160 199442 164212
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 202690 150396 202696 150408
rect 3384 150368 202696 150396
rect 3384 150356 3390 150368
rect 202690 150356 202696 150368
rect 202748 150356 202754 150408
rect 296070 139340 296076 139392
rect 296128 139380 296134 139392
rect 580166 139380 580172 139392
rect 296128 139352 580172 139380
rect 296128 139340 296134 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 266998 126896 267004 126948
rect 267056 126936 267062 126948
rect 580166 126936 580172 126948
rect 267056 126908 580172 126936
rect 267056 126896 267062 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 265710 113092 265716 113144
rect 265768 113132 265774 113144
rect 579798 113132 579804 113144
rect 265768 113104 579804 113132
rect 265768 113092 265774 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 200758 111772 200764 111784
rect 3200 111744 200764 111772
rect 3200 111732 3206 111744
rect 200758 111732 200764 111744
rect 200816 111732 200822 111784
rect 296162 100648 296168 100700
rect 296220 100688 296226 100700
rect 580166 100688 580172 100700
rect 296220 100660 580172 100688
rect 296220 100648 296226 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 202506 97968 202512 97980
rect 3292 97940 202512 97968
rect 3292 97928 3298 97940
rect 202506 97928 202512 97940
rect 202564 97928 202570 97980
rect 249058 88952 249064 89004
rect 249116 88992 249122 89004
rect 502334 88992 502340 89004
rect 249116 88964 502340 88992
rect 249116 88952 249122 88964
rect 502334 88952 502340 88964
rect 502392 88952 502398 89004
rect 235350 87728 235356 87780
rect 235408 87768 235414 87780
rect 316126 87768 316132 87780
rect 235408 87740 316132 87768
rect 235408 87728 235414 87740
rect 316126 87728 316132 87740
rect 316184 87728 316190 87780
rect 242250 87660 242256 87712
rect 242308 87700 242314 87712
rect 407114 87700 407120 87712
rect 242308 87672 407120 87700
rect 242308 87660 242314 87672
rect 407114 87660 407120 87672
rect 407172 87660 407178 87712
rect 244918 87592 244924 87644
rect 244976 87632 244982 87644
rect 448514 87632 448520 87644
rect 244976 87604 448520 87632
rect 244976 87592 244982 87604
rect 448514 87592 448520 87604
rect 448572 87592 448578 87644
rect 264238 86912 264244 86964
rect 264296 86952 264302 86964
rect 580166 86952 580172 86964
rect 264296 86924 580172 86952
rect 264296 86912 264302 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 247586 86300 247592 86352
rect 247644 86340 247650 86352
rect 481634 86340 481640 86352
rect 247644 86312 481640 86340
rect 247644 86300 247650 86312
rect 481634 86300 481640 86312
rect 481692 86300 481698 86352
rect 250346 86232 250352 86284
rect 250404 86272 250410 86284
rect 514846 86272 514852 86284
rect 250404 86244 514852 86272
rect 250404 86232 250410 86244
rect 514846 86232 514852 86244
rect 514904 86232 514910 86284
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 202414 85524 202420 85536
rect 3384 85496 202420 85524
rect 3384 85484 3390 85496
rect 202414 85484 202420 85496
rect 202472 85484 202478 85536
rect 239398 84872 239404 84924
rect 239456 84912 239462 84924
rect 285674 84912 285680 84924
rect 239456 84884 285680 84912
rect 239456 84872 239462 84884
rect 285674 84872 285680 84884
rect 285732 84872 285738 84924
rect 254486 84804 254492 84856
rect 254544 84844 254550 84856
rect 563054 84844 563060 84856
rect 254544 84816 563060 84844
rect 254544 84804 254550 84816
rect 563054 84804 563060 84816
rect 563112 84804 563118 84856
rect 242158 83444 242164 83496
rect 242216 83484 242222 83496
rect 402974 83484 402980 83496
rect 242216 83456 402980 83484
rect 242216 83444 242222 83456
rect 402974 83444 402980 83456
rect 403032 83444 403038 83496
rect 230934 82152 230940 82204
rect 230992 82192 230998 82204
rect 262214 82192 262220 82204
rect 230992 82164 262220 82192
rect 230992 82152 230998 82164
rect 262214 82152 262220 82164
rect 262272 82152 262278 82204
rect 247494 82084 247500 82136
rect 247552 82124 247558 82136
rect 477494 82124 477500 82136
rect 247552 82096 477500 82124
rect 247552 82084 247558 82096
rect 477494 82084 477500 82096
rect 477552 82084 477558 82136
rect 265618 73108 265624 73160
rect 265676 73148 265682 73160
rect 580166 73148 580172 73160
rect 265676 73120 580172 73148
rect 265676 73108 265682 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 202322 71720 202328 71732
rect 3384 71692 202328 71720
rect 3384 71680 3390 71692
rect 202322 71680 202328 71692
rect 202380 71680 202386 71732
rect 295978 60664 295984 60716
rect 296036 60704 296042 60716
rect 580166 60704 580172 60716
rect 296036 60676 580172 60704
rect 296036 60664 296042 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3326 59304 3332 59356
rect 3384 59344 3390 59356
rect 202230 59344 202236 59356
rect 3384 59316 202236 59344
rect 3384 59304 3390 59316
rect 202230 59304 202236 59316
rect 202288 59304 202294 59356
rect 202966 58624 202972 58676
rect 203024 58664 203030 58676
rect 580258 58664 580264 58676
rect 203024 58636 580264 58664
rect 203024 58624 203030 58636
rect 580258 58624 580264 58636
rect 580316 58624 580322 58676
rect 260098 48968 260104 49020
rect 260156 49008 260162 49020
rect 454034 49008 454040 49020
rect 260156 48980 454040 49008
rect 260156 48968 260162 48980
rect 454034 48968 454040 48980
rect 454092 48968 454098 49020
rect 211614 46248 211620 46300
rect 211672 46288 211678 46300
rect 226702 46288 226708 46300
rect 211672 46260 226708 46288
rect 211672 46248 211678 46260
rect 226702 46248 226708 46260
rect 226760 46248 226766 46300
rect 160094 46180 160100 46232
rect 160152 46220 160158 46232
rect 222654 46220 222660 46232
rect 160152 46192 222660 46220
rect 160152 46180 160158 46192
rect 222654 46180 222660 46192
rect 222712 46180 222718 46232
rect 124214 37884 124220 37936
rect 124272 37924 124278 37936
rect 208118 37924 208124 37936
rect 124272 37896 208124 37924
rect 124272 37884 124278 37896
rect 208118 37884 208124 37896
rect 208176 37884 208182 37936
rect 95234 35164 95240 35216
rect 95292 35204 95298 35216
rect 209130 35204 209136 35216
rect 95292 35176 209136 35204
rect 95292 35164 95298 35176
rect 209130 35164 209136 35176
rect 209188 35164 209194 35216
rect 258718 35164 258724 35216
rect 258776 35204 258782 35216
rect 442994 35204 443000 35216
rect 258776 35176 443000 35204
rect 258776 35164 258782 35176
rect 442994 35164 443000 35176
rect 443052 35164 443058 35216
rect 202874 33056 202880 33108
rect 202932 33096 202938 33108
rect 580166 33096 580172 33108
rect 202932 33068 580172 33096
rect 202932 33056 202938 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 203518 33028 203524 33040
rect 3476 33000 203524 33028
rect 3476 32988 3482 33000
rect 203518 32988 203524 33000
rect 203576 32988 203582 33040
rect 256234 28296 256240 28348
rect 256292 28336 256298 28348
rect 494054 28336 494060 28348
rect 256292 28308 494060 28336
rect 256292 28296 256298 28308
rect 494054 28296 494060 28308
rect 494112 28296 494118 28348
rect 248966 28228 248972 28280
rect 249024 28268 249030 28280
rect 498194 28268 498200 28280
rect 249024 28240 498200 28268
rect 249024 28228 249030 28240
rect 498194 28228 498200 28240
rect 498252 28228 498258 28280
rect 256142 26936 256148 26988
rect 256200 26976 256206 26988
rect 407206 26976 407212 26988
rect 256200 26948 407212 26976
rect 256200 26936 256206 26948
rect 407206 26936 407212 26948
rect 407264 26936 407270 26988
rect 256050 26868 256056 26920
rect 256108 26908 256114 26920
rect 415394 26908 415400 26920
rect 256108 26880 415400 26908
rect 256108 26868 256114 26880
rect 415394 26868 415400 26880
rect 415452 26868 415458 26920
rect 232498 25984 232504 26036
rect 232556 26024 232562 26036
rect 287054 26024 287060 26036
rect 232556 25996 287060 26024
rect 232556 25984 232562 25996
rect 287054 25984 287060 25996
rect 287112 25984 287118 26036
rect 235166 25916 235172 25968
rect 235224 25956 235230 25968
rect 311894 25956 311900 25968
rect 235224 25928 311900 25956
rect 235224 25916 235230 25928
rect 311894 25916 311900 25928
rect 311952 25916 311958 25968
rect 235074 25848 235080 25900
rect 235132 25888 235138 25900
rect 322934 25888 322940 25900
rect 235132 25860 322940 25888
rect 235132 25848 235138 25860
rect 322934 25848 322940 25860
rect 322992 25848 322998 25900
rect 236454 25780 236460 25832
rect 236512 25820 236518 25832
rect 332594 25820 332600 25832
rect 236512 25792 332600 25820
rect 236512 25780 236518 25792
rect 332594 25780 332600 25792
rect 332652 25780 332658 25832
rect 239122 25712 239128 25764
rect 239180 25752 239186 25764
rect 375374 25752 375380 25764
rect 239180 25724 375380 25752
rect 239180 25712 239186 25724
rect 375374 25712 375380 25724
rect 375432 25712 375438 25764
rect 243538 25644 243544 25696
rect 243596 25684 243602 25696
rect 425054 25684 425060 25696
rect 243596 25656 425060 25684
rect 243596 25644 243602 25656
rect 425054 25644 425060 25656
rect 425112 25644 425118 25696
rect 244734 25576 244740 25628
rect 244792 25616 244798 25628
rect 440234 25616 440240 25628
rect 244792 25588 440240 25616
rect 244792 25576 244798 25588
rect 440234 25576 440240 25588
rect 440292 25576 440298 25628
rect 244826 25508 244832 25560
rect 244884 25548 244890 25560
rect 447134 25548 447140 25560
rect 244884 25520 447140 25548
rect 244884 25508 244890 25520
rect 447134 25508 447140 25520
rect 447192 25508 447198 25560
rect 232406 24488 232412 24540
rect 232464 24528 232470 24540
rect 276014 24528 276020 24540
rect 232464 24500 276020 24528
rect 232464 24488 232470 24500
rect 276014 24488 276020 24500
rect 276072 24488 276078 24540
rect 232314 24420 232320 24472
rect 232372 24460 232378 24472
rect 280154 24460 280160 24472
rect 232372 24432 280160 24460
rect 232372 24420 232378 24432
rect 280154 24420 280160 24432
rect 280212 24420 280218 24472
rect 250254 24352 250260 24404
rect 250312 24392 250318 24404
rect 517514 24392 517520 24404
rect 250312 24364 517520 24392
rect 250312 24352 250318 24364
rect 517514 24352 517520 24364
rect 517572 24352 517578 24404
rect 253106 24284 253112 24336
rect 253164 24324 253170 24336
rect 542354 24324 542360 24336
rect 253164 24296 542360 24324
rect 253164 24284 253170 24296
rect 542354 24284 542360 24296
rect 542412 24284 542418 24336
rect 253198 24216 253204 24268
rect 253256 24256 253262 24268
rect 546494 24256 546500 24268
rect 253256 24228 546500 24256
rect 253256 24216 253262 24228
rect 546494 24216 546500 24228
rect 546552 24216 546558 24268
rect 253014 24148 253020 24200
rect 253072 24188 253078 24200
rect 553394 24188 553400 24200
rect 253072 24160 553400 24188
rect 253072 24148 253078 24160
rect 553394 24148 553400 24160
rect 553452 24148 553458 24200
rect 254394 24080 254400 24132
rect 254452 24120 254458 24132
rect 564526 24120 564532 24132
rect 254452 24092 564532 24120
rect 254452 24080 254458 24092
rect 564526 24080 564532 24092
rect 564584 24080 564590 24132
rect 236362 23128 236368 23180
rect 236420 23168 236426 23180
rect 336734 23168 336740 23180
rect 236420 23140 336740 23168
rect 236420 23128 236426 23140
rect 336734 23128 336740 23140
rect 336792 23128 336798 23180
rect 246114 23060 246120 23112
rect 246172 23100 246178 23112
rect 463694 23100 463700 23112
rect 246172 23072 463700 23100
rect 246172 23060 246178 23072
rect 463694 23060 463700 23072
rect 463752 23060 463758 23112
rect 247402 22992 247408 23044
rect 247460 23032 247466 23044
rect 473354 23032 473360 23044
rect 247460 23004 473360 23032
rect 247460 22992 247466 23004
rect 473354 22992 473360 23004
rect 473412 22992 473418 23044
rect 248782 22924 248788 22976
rect 248840 22964 248846 22976
rect 490006 22964 490012 22976
rect 248840 22936 490012 22964
rect 248840 22924 248846 22936
rect 490006 22924 490012 22936
rect 490064 22924 490070 22976
rect 248874 22856 248880 22908
rect 248932 22896 248938 22908
rect 496814 22896 496820 22908
rect 248932 22868 496820 22896
rect 248932 22856 248938 22868
rect 496814 22856 496820 22868
rect 496872 22856 496878 22908
rect 250162 22788 250168 22840
rect 250220 22828 250226 22840
rect 506566 22828 506572 22840
rect 250220 22800 506572 22828
rect 250220 22788 250226 22800
rect 506566 22788 506572 22800
rect 506624 22788 506630 22840
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 15838 22760 15844 22772
rect 5592 22732 15844 22760
rect 5592 22720 5598 22732
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 250070 22720 250076 22772
rect 250128 22760 250134 22772
rect 510614 22760 510620 22772
rect 250128 22732 510620 22760
rect 250128 22720 250134 22732
rect 510614 22720 510620 22732
rect 510672 22720 510678 22772
rect 241974 21836 241980 21888
rect 242032 21876 242038 21888
rect 409874 21876 409880 21888
rect 242032 21848 409880 21876
rect 242032 21836 242038 21848
rect 409874 21836 409880 21848
rect 409932 21836 409938 21888
rect 243446 21768 243452 21820
rect 243504 21808 243510 21820
rect 420914 21808 420920 21820
rect 243504 21780 420920 21808
rect 243504 21768 243510 21780
rect 420914 21768 420920 21780
rect 420972 21768 420978 21820
rect 243354 21700 243360 21752
rect 243412 21740 243418 21752
rect 423674 21740 423680 21752
rect 243412 21712 423680 21740
rect 243412 21700 243418 21712
rect 423674 21700 423680 21712
rect 423732 21700 423738 21752
rect 243262 21632 243268 21684
rect 243320 21672 243326 21684
rect 427814 21672 427820 21684
rect 243320 21644 427820 21672
rect 243320 21632 243326 21644
rect 427814 21632 427820 21644
rect 427872 21632 427878 21684
rect 244550 21564 244556 21616
rect 244608 21604 244614 21616
rect 438854 21604 438860 21616
rect 244608 21576 438860 21604
rect 244608 21564 244614 21576
rect 438854 21564 438860 21576
rect 438912 21564 438918 21616
rect 244642 21496 244648 21548
rect 244700 21536 244706 21548
rect 441614 21536 441620 21548
rect 244700 21508 441620 21536
rect 244700 21496 244706 21508
rect 441614 21496 441620 21508
rect 441672 21496 441678 21548
rect 246022 21428 246028 21480
rect 246080 21468 246086 21480
rect 456886 21468 456892 21480
rect 246080 21440 456892 21468
rect 246080 21428 246086 21440
rect 456886 21428 456892 21440
rect 456944 21428 456950 21480
rect 245930 21360 245936 21412
rect 245988 21400 245994 21412
rect 459554 21400 459560 21412
rect 245988 21372 459560 21400
rect 245988 21360 245994 21372
rect 459554 21360 459560 21372
rect 459612 21360 459618 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 202138 20652 202144 20664
rect 3476 20624 202144 20652
rect 3476 20612 3482 20624
rect 202138 20612 202144 20624
rect 202196 20612 202202 20664
rect 237742 20204 237748 20256
rect 237800 20244 237806 20256
rect 349246 20244 349252 20256
rect 237800 20216 349252 20244
rect 237800 20204 237806 20216
rect 349246 20204 349252 20216
rect 349304 20204 349310 20256
rect 237834 20136 237840 20188
rect 237892 20176 237898 20188
rect 353294 20176 353300 20188
rect 237892 20148 353300 20176
rect 237892 20136 237898 20148
rect 353294 20136 353300 20148
rect 353352 20136 353358 20188
rect 239030 20068 239036 20120
rect 239088 20108 239094 20120
rect 373994 20108 374000 20120
rect 239088 20080 374000 20108
rect 239088 20068 239094 20080
rect 373994 20068 374000 20080
rect 374052 20068 374058 20120
rect 240502 20000 240508 20052
rect 240560 20040 240566 20052
rect 389174 20040 389180 20052
rect 240560 20012 389180 20040
rect 240560 20000 240566 20012
rect 389174 20000 389180 20012
rect 389232 20000 389238 20052
rect 240410 19932 240416 19984
rect 240468 19972 240474 19984
rect 391934 19972 391940 19984
rect 240468 19944 391940 19972
rect 240468 19932 240474 19944
rect 391934 19932 391940 19944
rect 391992 19932 391998 19984
rect 233694 19048 233700 19100
rect 233752 19088 233758 19100
rect 296714 19088 296720 19100
rect 233752 19060 296720 19088
rect 233752 19048 233758 19060
rect 296714 19048 296720 19060
rect 296772 19048 296778 19100
rect 233602 18980 233608 19032
rect 233660 19020 233666 19032
rect 299474 19020 299480 19032
rect 233660 18992 299480 19020
rect 233660 18980 233666 18992
rect 299474 18980 299480 18992
rect 299532 18980 299538 19032
rect 233510 18912 233516 18964
rect 233568 18952 233574 18964
rect 303614 18952 303620 18964
rect 233568 18924 303620 18952
rect 233568 18912 233574 18924
rect 303614 18912 303620 18924
rect 303672 18912 303678 18964
rect 234798 18844 234804 18896
rect 234856 18884 234862 18896
rect 314654 18884 314660 18896
rect 234856 18856 314660 18884
rect 234856 18844 234862 18856
rect 314654 18844 314660 18856
rect 314712 18844 314718 18896
rect 234982 18776 234988 18828
rect 235040 18816 235046 18828
rect 317414 18816 317420 18828
rect 235040 18788 317420 18816
rect 235040 18776 235046 18788
rect 317414 18776 317420 18788
rect 317472 18776 317478 18828
rect 234890 18708 234896 18760
rect 234948 18748 234954 18760
rect 321554 18748 321560 18760
rect 234948 18720 321560 18748
rect 234948 18708 234954 18720
rect 321554 18708 321560 18720
rect 321612 18708 321618 18760
rect 236178 18640 236184 18692
rect 236236 18680 236242 18692
rect 332686 18680 332692 18692
rect 236236 18652 332692 18680
rect 236236 18640 236242 18652
rect 332686 18640 332692 18652
rect 332744 18640 332750 18692
rect 236270 18572 236276 18624
rect 236328 18612 236334 18624
rect 335354 18612 335360 18624
rect 236328 18584 335360 18612
rect 236328 18572 236334 18584
rect 335354 18572 335360 18584
rect 335412 18572 335418 18624
rect 232130 17620 232136 17672
rect 232188 17660 232194 17672
rect 278774 17660 278780 17672
rect 232188 17632 278780 17660
rect 232188 17620 232194 17632
rect 278774 17620 278780 17632
rect 278832 17620 278838 17672
rect 232222 17552 232228 17604
rect 232280 17592 232286 17604
rect 282914 17592 282920 17604
rect 232280 17564 282920 17592
rect 232280 17552 232286 17564
rect 282914 17552 282920 17564
rect 282972 17552 282978 17604
rect 251542 17484 251548 17536
rect 251600 17524 251606 17536
rect 534074 17524 534080 17536
rect 251600 17496 534080 17524
rect 251600 17484 251606 17496
rect 534074 17484 534080 17496
rect 534132 17484 534138 17536
rect 252738 17416 252744 17468
rect 252796 17456 252802 17468
rect 545114 17456 545120 17468
rect 252796 17428 545120 17456
rect 252796 17416 252802 17428
rect 545114 17416 545120 17428
rect 545172 17416 545178 17468
rect 252922 17348 252928 17400
rect 252980 17388 252986 17400
rect 547874 17388 547880 17400
rect 252980 17360 547880 17388
rect 252980 17348 252986 17360
rect 547874 17348 547880 17360
rect 547932 17348 547938 17400
rect 252830 17280 252836 17332
rect 252888 17320 252894 17332
rect 552014 17320 552020 17332
rect 252888 17292 552020 17320
rect 252888 17280 252894 17292
rect 552014 17280 552020 17292
rect 552072 17280 552078 17332
rect 180794 17212 180800 17264
rect 180852 17252 180858 17264
rect 224034 17252 224040 17264
rect 180852 17224 224040 17252
rect 180852 17212 180858 17224
rect 224034 17212 224040 17224
rect 224092 17212 224098 17264
rect 254302 17212 254308 17264
rect 254360 17252 254366 17264
rect 567194 17252 567200 17264
rect 254360 17224 567200 17252
rect 254360 17212 254366 17224
rect 567194 17212 567200 17224
rect 567252 17212 567258 17264
rect 243170 16260 243176 16312
rect 243228 16300 243234 16312
rect 418522 16300 418528 16312
rect 243228 16272 418528 16300
rect 243228 16260 243234 16272
rect 418522 16260 418528 16272
rect 418580 16260 418586 16312
rect 248690 16192 248696 16244
rect 248748 16232 248754 16244
rect 498930 16232 498936 16244
rect 248748 16204 498936 16232
rect 248748 16192 248754 16204
rect 498930 16192 498936 16204
rect 498988 16192 498994 16244
rect 249886 16124 249892 16176
rect 249944 16164 249950 16176
rect 509602 16164 509608 16176
rect 249944 16136 509608 16164
rect 249944 16124 249950 16136
rect 509602 16124 509608 16136
rect 509660 16124 509666 16176
rect 136450 16056 136456 16108
rect 136508 16096 136514 16108
rect 220170 16096 220176 16108
rect 136508 16068 220176 16096
rect 136508 16056 136514 16068
rect 220170 16056 220176 16068
rect 220228 16056 220234 16108
rect 249794 16056 249800 16108
rect 249852 16096 249858 16108
rect 513374 16096 513380 16108
rect 249852 16068 513380 16096
rect 249852 16056 249858 16068
rect 513374 16056 513380 16068
rect 513432 16056 513438 16108
rect 71498 15988 71504 16040
rect 71556 16028 71562 16040
rect 210510 16028 210516 16040
rect 71556 16000 210516 16028
rect 71556 15988 71562 16000
rect 210510 15988 210516 16000
rect 210568 15988 210574 16040
rect 249978 15988 249984 16040
rect 250036 16028 250042 16040
rect 517146 16028 517152 16040
rect 250036 16000 517152 16028
rect 250036 15988 250042 16000
rect 517146 15988 517152 16000
rect 517204 15988 517210 16040
rect 35986 15920 35992 15972
rect 36044 15960 36050 15972
rect 212810 15960 212816 15972
rect 36044 15932 212816 15960
rect 36044 15920 36050 15932
rect 212810 15920 212816 15932
rect 212868 15920 212874 15972
rect 251450 15920 251456 15972
rect 251508 15960 251514 15972
rect 527818 15960 527824 15972
rect 251508 15932 527824 15960
rect 251508 15920 251514 15932
rect 527818 15920 527824 15932
rect 527876 15920 527882 15972
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 210234 15892 210240 15904
rect 9732 15864 210240 15892
rect 9732 15852 9738 15864
rect 210234 15852 210240 15864
rect 210292 15852 210298 15904
rect 251358 15852 251364 15904
rect 251416 15892 251422 15904
rect 531406 15892 531412 15904
rect 251416 15864 531412 15892
rect 251416 15852 251422 15864
rect 531406 15852 531412 15864
rect 531464 15852 531470 15904
rect 163498 14968 163504 15020
rect 163556 15008 163562 15020
rect 218422 15008 218428 15020
rect 163556 14980 218428 15008
rect 163556 14968 163562 14980
rect 218422 14968 218428 14980
rect 218480 14968 218486 15020
rect 112346 14900 112352 14952
rect 112404 14940 112410 14952
rect 218514 14940 218520 14952
rect 112404 14912 218520 14940
rect 112404 14900 112410 14912
rect 218514 14900 218520 14912
rect 218572 14900 218578 14952
rect 98178 14832 98184 14884
rect 98236 14872 98242 14884
rect 217226 14872 217232 14884
rect 98236 14844 217232 14872
rect 98236 14832 98242 14844
rect 217226 14832 217232 14844
rect 217284 14832 217290 14884
rect 91554 14764 91560 14816
rect 91612 14804 91618 14816
rect 217134 14804 217140 14816
rect 91612 14776 217140 14804
rect 91612 14764 91618 14776
rect 217134 14764 217140 14776
rect 217192 14764 217198 14816
rect 247126 14764 247132 14816
rect 247184 14804 247190 14816
rect 473446 14804 473452 14816
rect 247184 14776 473452 14804
rect 247184 14764 247190 14776
rect 473446 14764 473452 14776
rect 473504 14764 473510 14816
rect 74994 14696 75000 14748
rect 75052 14736 75058 14748
rect 215662 14736 215668 14748
rect 75052 14708 215668 14736
rect 75052 14696 75058 14708
rect 215662 14696 215668 14708
rect 215720 14696 215726 14748
rect 247218 14696 247224 14748
rect 247276 14736 247282 14748
rect 476482 14736 476488 14748
rect 247276 14708 476488 14736
rect 247276 14696 247282 14708
rect 476482 14696 476488 14708
rect 476540 14696 476546 14748
rect 44174 14628 44180 14680
rect 44232 14668 44238 14680
rect 211798 14668 211804 14680
rect 44232 14640 211804 14668
rect 44232 14628 44238 14640
rect 211798 14628 211804 14640
rect 211856 14628 211862 14680
rect 247310 14628 247316 14680
rect 247368 14668 247374 14680
rect 481726 14668 481732 14680
rect 247368 14640 481732 14668
rect 247368 14628 247374 14640
rect 481726 14628 481732 14640
rect 481784 14628 481790 14680
rect 27706 14560 27712 14612
rect 27764 14600 27770 14612
rect 211430 14600 211436 14612
rect 27764 14572 211436 14600
rect 27764 14560 27770 14572
rect 211430 14560 211436 14572
rect 211488 14560 211494 14612
rect 248506 14560 248512 14612
rect 248564 14600 248570 14612
rect 492306 14600 492312 14612
rect 248564 14572 492312 14600
rect 248564 14560 248570 14572
rect 492306 14560 492312 14572
rect 492364 14560 492370 14612
rect 22554 14492 22560 14544
rect 22612 14532 22618 14544
rect 211338 14532 211344 14544
rect 22612 14504 211344 14532
rect 22612 14492 22618 14504
rect 211338 14492 211344 14504
rect 211396 14492 211402 14544
rect 248598 14492 248604 14544
rect 248656 14532 248662 14544
rect 495434 14532 495440 14544
rect 248656 14504 495440 14532
rect 248656 14492 248662 14504
rect 495434 14492 495440 14504
rect 495492 14492 495498 14544
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 211522 14464 211528 14476
rect 18012 14436 211528 14464
rect 18012 14424 18018 14436
rect 211522 14424 211528 14436
rect 211580 14424 211586 14476
rect 254210 14424 254216 14476
rect 254268 14464 254274 14476
rect 570322 14464 570328 14476
rect 254268 14436 570328 14464
rect 254268 14424 254274 14436
rect 570322 14424 570328 14436
rect 570380 14424 570386 14476
rect 80882 13472 80888 13524
rect 80940 13512 80946 13524
rect 215570 13512 215576 13524
rect 80940 13484 215576 13512
rect 80940 13472 80946 13484
rect 215570 13472 215576 13484
rect 215628 13472 215634 13524
rect 243078 13472 243084 13524
rect 243136 13512 243142 13524
rect 430850 13512 430856 13524
rect 243136 13484 430856 13512
rect 243136 13472 243142 13484
rect 430850 13472 430856 13484
rect 430908 13472 430914 13524
rect 63218 13404 63224 13456
rect 63276 13444 63282 13456
rect 214374 13444 214380 13456
rect 63276 13416 214380 13444
rect 63276 13404 63282 13416
rect 214374 13404 214380 13416
rect 214432 13404 214438 13456
rect 244274 13404 244280 13456
rect 244332 13444 244338 13456
rect 440326 13444 440332 13456
rect 244332 13416 440332 13444
rect 244332 13404 244338 13416
rect 440326 13404 440332 13416
rect 440384 13404 440390 13456
rect 59354 13336 59360 13388
rect 59412 13376 59418 13388
rect 214466 13376 214472 13388
rect 59412 13348 214472 13376
rect 59412 13336 59418 13348
rect 214466 13336 214472 13348
rect 214524 13336 214530 13388
rect 244458 13336 244464 13388
rect 244516 13376 244522 13388
rect 445018 13376 445024 13388
rect 244516 13348 445024 13376
rect 244516 13336 244522 13348
rect 445018 13336 445024 13348
rect 445076 13336 445082 13388
rect 56042 13268 56048 13320
rect 56100 13308 56106 13320
rect 214558 13308 214564 13320
rect 56100 13280 214564 13308
rect 56100 13268 56106 13280
rect 214558 13268 214564 13280
rect 214616 13268 214622 13320
rect 244366 13268 244372 13320
rect 244424 13308 244430 13320
rect 448606 13308 448612 13320
rect 244424 13280 448612 13308
rect 244424 13268 244430 13280
rect 448606 13268 448612 13280
rect 448664 13268 448670 13320
rect 52546 13200 52552 13252
rect 52604 13240 52610 13252
rect 214282 13240 214288 13252
rect 52604 13212 214288 13240
rect 52604 13200 52610 13212
rect 214282 13200 214288 13212
rect 214340 13200 214346 13252
rect 245746 13200 245752 13252
rect 245804 13240 245810 13252
rect 459186 13240 459192 13252
rect 245804 13212 459192 13240
rect 245804 13200 245810 13212
rect 459186 13200 459192 13212
rect 459244 13200 459250 13252
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 210050 13172 210056 13184
rect 8812 13144 210056 13172
rect 8812 13132 8818 13144
rect 210050 13132 210056 13144
rect 210108 13132 210114 13184
rect 245654 13132 245660 13184
rect 245712 13172 245718 13184
rect 462314 13172 462320 13184
rect 245712 13144 462320 13172
rect 245712 13132 245718 13144
rect 462314 13132 462320 13144
rect 462372 13132 462378 13184
rect 3418 13064 3424 13116
rect 3476 13104 3482 13116
rect 210142 13104 210148 13116
rect 3476 13076 210148 13104
rect 3476 13064 3482 13076
rect 210142 13064 210148 13076
rect 210200 13064 210206 13116
rect 245838 13064 245844 13116
rect 245896 13104 245902 13116
rect 465810 13104 465816 13116
rect 245896 13076 465816 13104
rect 245896 13064 245902 13076
rect 465810 13064 465816 13076
rect 465868 13064 465874 13116
rect 114738 12180 114744 12232
rect 114796 12220 114802 12232
rect 218238 12220 218244 12232
rect 114796 12192 218244 12220
rect 114796 12180 114802 12192
rect 218238 12180 218244 12192
rect 218296 12180 218302 12232
rect 110414 12112 110420 12164
rect 110472 12152 110478 12164
rect 218330 12152 218336 12164
rect 110472 12124 218336 12152
rect 110472 12112 110478 12124
rect 218330 12112 218336 12124
rect 218388 12112 218394 12164
rect 108114 12044 108120 12096
rect 108172 12084 108178 12096
rect 218882 12084 218888 12096
rect 108172 12056 218888 12084
rect 108172 12044 108178 12056
rect 218882 12044 218888 12056
rect 218940 12044 218946 12096
rect 240318 12044 240324 12096
rect 240376 12084 240382 12096
rect 395338 12084 395344 12096
rect 240376 12056 395344 12084
rect 240376 12044 240382 12056
rect 395338 12044 395344 12056
rect 395396 12044 395402 12096
rect 44266 11976 44272 12028
rect 44324 12016 44330 12028
rect 212718 12016 212724 12028
rect 44324 11988 212724 12016
rect 44324 11976 44330 11988
rect 212718 11976 212724 11988
rect 212776 11976 212782 12028
rect 241698 11976 241704 12028
rect 241756 12016 241762 12028
rect 402514 12016 402520 12028
rect 241756 11988 402520 12016
rect 241756 11976 241762 11988
rect 402514 11976 402520 11988
rect 402572 11976 402578 12028
rect 36722 11908 36728 11960
rect 36780 11948 36786 11960
rect 213086 11948 213092 11960
rect 36780 11920 213092 11948
rect 36780 11908 36786 11920
rect 213086 11908 213092 11920
rect 213144 11908 213150 11960
rect 241882 11908 241888 11960
rect 241940 11948 241946 11960
rect 406010 11948 406016 11960
rect 241940 11920 406016 11948
rect 241940 11908 241946 11920
rect 406010 11908 406016 11920
rect 406068 11908 406074 11960
rect 33594 11840 33600 11892
rect 33652 11880 33658 11892
rect 213454 11880 213460 11892
rect 33652 11852 213460 11880
rect 33652 11840 33658 11852
rect 213454 11840 213460 11852
rect 213512 11840 213518 11892
rect 241790 11840 241796 11892
rect 241848 11880 241854 11892
rect 409138 11880 409144 11892
rect 241848 11852 409144 11880
rect 241848 11840 241854 11852
rect 409138 11840 409144 11852
rect 409196 11840 409202 11892
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 212350 11812 212356 11824
rect 26292 11784 212356 11812
rect 26292 11772 26298 11784
rect 212350 11772 212356 11784
rect 212408 11772 212414 11824
rect 242986 11772 242992 11824
rect 243044 11812 243050 11824
rect 423766 11812 423772 11824
rect 243044 11784 423772 11812
rect 243044 11772 243050 11784
rect 423766 11772 423772 11784
rect 423824 11772 423830 11824
rect 21818 11704 21824 11756
rect 21876 11744 21882 11756
rect 211246 11744 211252 11756
rect 21876 11716 211252 11744
rect 21876 11704 21882 11716
rect 211246 11704 211252 11716
rect 211304 11704 211310 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 426802 11744 426808 11756
rect 242952 11716 426808 11744
rect 242952 11704 242958 11716
rect 426802 11704 426808 11716
rect 426860 11704 426866 11756
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 159358 10752 159364 10804
rect 159416 10792 159422 10804
rect 218790 10792 218796 10804
rect 159416 10764 218796 10792
rect 159416 10752 159422 10764
rect 218790 10752 218796 10764
rect 218848 10752 218854 10804
rect 97442 10684 97448 10736
rect 97500 10724 97506 10736
rect 216858 10724 216864 10736
rect 97500 10696 216864 10724
rect 97500 10684 97506 10696
rect 216858 10684 216864 10696
rect 216916 10684 216922 10736
rect 93946 10616 93952 10668
rect 94004 10656 94010 10668
rect 217042 10656 217048 10668
rect 94004 10628 217048 10656
rect 94004 10616 94010 10628
rect 217042 10616 217048 10628
rect 217100 10616 217106 10668
rect 238938 10616 238944 10668
rect 238996 10656 239002 10668
rect 365806 10656 365812 10668
rect 238996 10628 365812 10656
rect 238996 10616 239002 10628
rect 365806 10616 365812 10628
rect 365864 10616 365870 10668
rect 89898 10548 89904 10600
rect 89956 10588 89962 10600
rect 216950 10588 216956 10600
rect 89956 10560 216956 10588
rect 89956 10548 89962 10560
rect 216950 10548 216956 10560
rect 217008 10548 217014 10600
rect 238846 10548 238852 10600
rect 238904 10588 238910 10600
rect 370130 10588 370136 10600
rect 238904 10560 370136 10588
rect 238904 10548 238910 10560
rect 370130 10548 370136 10560
rect 370188 10548 370194 10600
rect 86402 10480 86408 10532
rect 86460 10520 86466 10532
rect 216766 10520 216772 10532
rect 86460 10492 216772 10520
rect 86460 10480 86466 10492
rect 216766 10480 216772 10492
rect 216824 10480 216830 10532
rect 238754 10480 238760 10532
rect 238812 10520 238818 10532
rect 374086 10520 374092 10532
rect 238812 10492 374092 10520
rect 238812 10480 238818 10492
rect 374086 10480 374092 10492
rect 374144 10480 374150 10532
rect 75914 10412 75920 10464
rect 75972 10452 75978 10464
rect 216122 10452 216128 10464
rect 75972 10424 216128 10452
rect 75972 10412 75978 10424
rect 216122 10412 216128 10424
rect 216180 10412 216186 10464
rect 240134 10412 240140 10464
rect 240192 10452 240198 10464
rect 387794 10452 387800 10464
rect 240192 10424 387800 10452
rect 240192 10412 240198 10424
rect 387794 10412 387800 10424
rect 387852 10412 387858 10464
rect 72602 10344 72608 10396
rect 72660 10384 72666 10396
rect 215478 10384 215484 10396
rect 72660 10356 215484 10384
rect 72660 10344 72666 10356
rect 215478 10344 215484 10356
rect 215536 10344 215542 10396
rect 240226 10344 240232 10396
rect 240284 10384 240290 10396
rect 390646 10384 390652 10396
rect 240284 10356 390652 10384
rect 240284 10344 240290 10356
rect 390646 10344 390652 10356
rect 390704 10344 390710 10396
rect 69106 10276 69112 10328
rect 69164 10316 69170 10328
rect 215386 10316 215392 10328
rect 69164 10288 215392 10316
rect 69164 10276 69170 10288
rect 215386 10276 215392 10288
rect 215444 10276 215450 10328
rect 255498 10276 255504 10328
rect 255556 10316 255562 10328
rect 581730 10316 581736 10328
rect 255556 10288 581736 10316
rect 255556 10276 255562 10288
rect 581730 10276 581736 10288
rect 581788 10276 581794 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 156506 9392 156512 9444
rect 156564 9432 156570 9444
rect 222562 9432 222568 9444
rect 156564 9404 222568 9432
rect 156564 9392 156570 9404
rect 222562 9392 222568 9404
rect 222620 9392 222626 9444
rect 234706 9392 234712 9444
rect 234764 9432 234770 9444
rect 320910 9432 320916 9444
rect 234764 9404 320916 9432
rect 234764 9392 234770 9404
rect 320910 9392 320916 9404
rect 320968 9392 320974 9444
rect 149514 9324 149520 9376
rect 149572 9364 149578 9376
rect 221274 9364 221280 9376
rect 149572 9336 221280 9364
rect 149572 9324 149578 9336
rect 221274 9324 221280 9336
rect 221332 9324 221338 9376
rect 236086 9324 236092 9376
rect 236144 9364 236150 9376
rect 338666 9364 338672 9376
rect 236144 9336 338672 9364
rect 236144 9324 236150 9336
rect 338666 9324 338672 9336
rect 338724 9324 338730 9376
rect 142430 9256 142436 9308
rect 142488 9296 142494 9308
rect 221182 9296 221188 9308
rect 142488 9268 221188 9296
rect 142488 9256 142494 9268
rect 221182 9256 221188 9268
rect 221240 9256 221246 9308
rect 235994 9256 236000 9308
rect 236052 9296 236058 9308
rect 342162 9296 342168 9308
rect 236052 9268 342168 9296
rect 236052 9256 236058 9268
rect 342162 9256 342168 9268
rect 342220 9256 342226 9308
rect 62022 9188 62028 9240
rect 62080 9228 62086 9240
rect 214190 9228 214196 9240
rect 62080 9200 214196 9228
rect 62080 9188 62086 9200
rect 214190 9188 214196 9200
rect 214248 9188 214254 9240
rect 237650 9188 237656 9240
rect 237708 9228 237714 9240
rect 352834 9228 352840 9240
rect 237708 9200 352840 9228
rect 237708 9188 237714 9200
rect 352834 9188 352840 9200
rect 352892 9188 352898 9240
rect 54938 9120 54944 9172
rect 54996 9160 55002 9172
rect 214098 9160 214104 9172
rect 54996 9132 214104 9160
rect 54996 9120 55002 9132
rect 214098 9120 214104 9132
rect 214156 9120 214162 9172
rect 237466 9120 237472 9172
rect 237524 9160 237530 9172
rect 356330 9160 356336 9172
rect 237524 9132 356336 9160
rect 237524 9120 237530 9132
rect 356330 9120 356336 9132
rect 356388 9120 356394 9172
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 210786 9092 210792 9104
rect 7708 9064 210792 9092
rect 7708 9052 7714 9064
rect 210786 9052 210792 9064
rect 210844 9052 210850 9104
rect 237558 9052 237564 9104
rect 237616 9092 237622 9104
rect 359918 9092 359924 9104
rect 237616 9064 359924 9092
rect 237616 9052 237622 9064
rect 359918 9052 359924 9064
rect 359976 9052 359982 9104
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 209958 9024 209964 9036
rect 2924 8996 209964 9024
rect 2924 8984 2930 8996
rect 209958 8984 209964 8996
rect 210016 8984 210022 9036
rect 261478 8984 261484 9036
rect 261536 9024 261542 9036
rect 475746 9024 475752 9036
rect 261536 8996 475752 9024
rect 261536 8984 261542 8996
rect 475746 8984 475752 8996
rect 475804 8984 475810 9036
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 209866 8956 209872 8968
rect 1728 8928 209872 8956
rect 1728 8916 1734 8928
rect 209866 8916 209872 8928
rect 209924 8916 209930 8968
rect 254118 8916 254124 8968
rect 254176 8956 254182 8968
rect 566826 8956 566832 8968
rect 254176 8928 566832 8956
rect 254176 8916 254182 8928
rect 566826 8916 566832 8928
rect 566884 8916 566890 8968
rect 202690 7964 202696 8016
rect 202748 8004 202754 8016
rect 225230 8004 225236 8016
rect 202748 7976 225236 8004
rect 202748 7964 202754 7976
rect 225230 7964 225236 7976
rect 225288 7964 225294 8016
rect 195606 7896 195612 7948
rect 195664 7936 195670 7948
rect 225322 7936 225328 7948
rect 195664 7908 225328 7936
rect 195664 7896 195670 7908
rect 225322 7896 225328 7908
rect 225380 7896 225386 7948
rect 167178 7828 167184 7880
rect 167236 7868 167242 7880
rect 222470 7868 222476 7880
rect 167236 7840 222476 7868
rect 167236 7828 167242 7840
rect 222470 7828 222476 7840
rect 222528 7828 222534 7880
rect 230842 7828 230848 7880
rect 230900 7868 230906 7880
rect 268838 7868 268844 7880
rect 230900 7840 268844 7868
rect 230900 7828 230906 7840
rect 268838 7828 268844 7840
rect 268896 7828 268902 7880
rect 158898 7760 158904 7812
rect 158956 7800 158962 7812
rect 222378 7800 222384 7812
rect 158956 7772 222384 7800
rect 158956 7760 158962 7772
rect 222378 7760 222384 7772
rect 222436 7760 222442 7812
rect 232038 7760 232044 7812
rect 232096 7800 232102 7812
rect 288986 7800 288992 7812
rect 232096 7772 288992 7800
rect 232096 7760 232102 7772
rect 288986 7760 288992 7772
rect 289044 7760 289050 7812
rect 148318 7692 148324 7744
rect 148376 7732 148382 7744
rect 220998 7732 221004 7744
rect 148376 7704 221004 7732
rect 148376 7692 148382 7704
rect 220998 7692 221004 7704
rect 221056 7692 221062 7744
rect 233326 7692 233332 7744
rect 233384 7732 233390 7744
rect 303154 7732 303160 7744
rect 233384 7704 303160 7732
rect 233384 7692 233390 7704
rect 303154 7692 303160 7704
rect 303212 7692 303218 7744
rect 144730 7624 144736 7676
rect 144788 7664 144794 7676
rect 221090 7664 221096 7676
rect 144788 7636 221096 7664
rect 144788 7624 144794 7636
rect 221090 7624 221096 7636
rect 221148 7624 221154 7676
rect 257430 7624 257436 7676
rect 257488 7664 257494 7676
rect 422570 7664 422576 7676
rect 257488 7636 422576 7664
rect 257488 7624 257494 7636
rect 422570 7624 422576 7636
rect 422628 7624 422634 7676
rect 121086 7556 121092 7608
rect 121144 7596 121150 7608
rect 217318 7596 217324 7608
rect 121144 7568 217324 7596
rect 121144 7556 121150 7568
rect 217318 7556 217324 7568
rect 217376 7556 217382 7608
rect 257522 7556 257528 7608
rect 257580 7596 257586 7608
rect 429654 7596 429660 7608
rect 257580 7568 429660 7596
rect 257580 7556 257586 7568
rect 429654 7556 429660 7568
rect 429712 7556 429718 7608
rect 230750 6672 230756 6724
rect 230808 6712 230814 6724
rect 265342 6712 265348 6724
rect 230808 6684 265348 6712
rect 230808 6672 230814 6684
rect 265342 6672 265348 6684
rect 265400 6672 265406 6724
rect 187326 6604 187332 6656
rect 187384 6644 187390 6656
rect 223758 6644 223764 6656
rect 187384 6616 223764 6644
rect 187384 6604 187390 6616
rect 223758 6604 223764 6616
rect 223816 6604 223822 6656
rect 230566 6604 230572 6656
rect 230624 6644 230630 6656
rect 267734 6644 267740 6656
rect 230624 6616 267740 6644
rect 230624 6604 230630 6616
rect 267734 6604 267740 6616
rect 267792 6604 267798 6656
rect 183738 6536 183744 6588
rect 183796 6576 183802 6588
rect 224402 6576 224408 6588
rect 183796 6548 224408 6576
rect 183796 6536 183802 6548
rect 224402 6536 224408 6548
rect 224460 6536 224466 6588
rect 230658 6536 230664 6588
rect 230716 6576 230722 6588
rect 271230 6576 271236 6588
rect 230716 6548 271236 6576
rect 230716 6536 230722 6548
rect 271230 6536 271236 6548
rect 271288 6536 271294 6588
rect 180242 6468 180248 6520
rect 180300 6508 180306 6520
rect 223850 6508 223856 6520
rect 180300 6480 223856 6508
rect 180300 6468 180306 6480
rect 223850 6468 223856 6480
rect 223908 6468 223914 6520
rect 231854 6468 231860 6520
rect 231912 6508 231918 6520
rect 285398 6508 285404 6520
rect 231912 6480 285404 6508
rect 231912 6468 231918 6480
rect 285398 6468 285404 6480
rect 285456 6468 285462 6520
rect 176654 6400 176660 6452
rect 176712 6440 176718 6452
rect 223942 6440 223948 6452
rect 176712 6412 223948 6440
rect 176712 6400 176718 6412
rect 223942 6400 223948 6412
rect 224000 6400 224006 6452
rect 241514 6400 241520 6452
rect 241572 6440 241578 6452
rect 404814 6440 404820 6452
rect 241572 6412 404820 6440
rect 241572 6400 241578 6412
rect 404814 6400 404820 6412
rect 404872 6400 404878 6452
rect 130562 6332 130568 6384
rect 130620 6372 130626 6384
rect 219802 6372 219808 6384
rect 130620 6344 219808 6372
rect 130620 6332 130626 6344
rect 219802 6332 219808 6344
rect 219860 6332 219866 6384
rect 241606 6332 241612 6384
rect 241664 6372 241670 6384
rect 411898 6372 411904 6384
rect 241664 6344 411904 6372
rect 241664 6332 241670 6344
rect 411898 6332 411904 6344
rect 411956 6332 411962 6384
rect 117590 6264 117596 6316
rect 117648 6304 117654 6316
rect 208026 6304 208032 6316
rect 117648 6276 208032 6304
rect 117648 6264 117654 6276
rect 208026 6264 208032 6276
rect 208084 6264 208090 6316
rect 231946 6264 231952 6316
rect 232004 6304 232010 6316
rect 281902 6304 281908 6316
rect 232004 6276 281908 6304
rect 232004 6264 232010 6276
rect 281902 6264 281908 6276
rect 281960 6264 281966 6316
rect 282178 6264 282184 6316
rect 282236 6304 282242 6316
rect 580994 6304 581000 6316
rect 282236 6276 581000 6304
rect 282236 6264 282242 6276
rect 580994 6264 581000 6276
rect 581052 6264 581058 6316
rect 92750 6196 92756 6248
rect 92808 6236 92814 6248
rect 217502 6236 217508 6248
rect 92808 6208 217508 6236
rect 92808 6196 92814 6208
rect 217502 6196 217508 6208
rect 217560 6196 217566 6248
rect 253934 6196 253940 6248
rect 253992 6236 253998 6248
rect 569126 6236 569132 6248
rect 253992 6208 569132 6236
rect 253992 6196 253998 6208
rect 569126 6196 569132 6208
rect 569184 6196 569190 6248
rect 25314 6128 25320 6180
rect 25372 6168 25378 6180
rect 188338 6168 188344 6180
rect 25372 6140 188344 6168
rect 25372 6128 25378 6140
rect 188338 6128 188344 6140
rect 188396 6128 188402 6180
rect 197906 6128 197912 6180
rect 197964 6168 197970 6180
rect 225138 6168 225144 6180
rect 197964 6140 225144 6168
rect 197964 6128 197970 6140
rect 225138 6128 225144 6140
rect 225196 6128 225202 6180
rect 254026 6128 254032 6180
rect 254084 6168 254090 6180
rect 572714 6168 572720 6180
rect 254084 6140 572720 6168
rect 254084 6128 254090 6140
rect 572714 6128 572720 6140
rect 572772 6128 572778 6180
rect 201402 5380 201408 5432
rect 201460 5420 201466 5432
rect 223482 5420 223488 5432
rect 201460 5392 223488 5420
rect 201460 5380 201466 5392
rect 223482 5380 223488 5392
rect 223540 5380 223546 5432
rect 187694 5312 187700 5364
rect 187752 5352 187758 5364
rect 219618 5352 219624 5364
rect 187752 5324 219624 5352
rect 187752 5312 187758 5324
rect 219618 5312 219624 5324
rect 219676 5312 219682 5364
rect 162486 5244 162492 5296
rect 162544 5284 162550 5296
rect 222930 5284 222936 5296
rect 162544 5256 222936 5284
rect 162544 5244 162550 5256
rect 222930 5244 222936 5256
rect 222988 5244 222994 5296
rect 150618 5176 150624 5228
rect 150676 5216 150682 5228
rect 220906 5216 220912 5228
rect 150676 5188 220912 5216
rect 150676 5176 150682 5188
rect 220906 5176 220912 5188
rect 220964 5176 220970 5228
rect 147122 5108 147128 5160
rect 147180 5148 147186 5160
rect 221550 5148 221556 5160
rect 147180 5120 221556 5148
rect 147180 5108 147186 5120
rect 221550 5108 221556 5120
rect 221608 5108 221614 5160
rect 237374 5108 237380 5160
rect 237432 5148 237438 5160
rect 355226 5148 355232 5160
rect 237432 5120 355232 5148
rect 237432 5108 237438 5120
rect 355226 5108 355232 5120
rect 355284 5108 355290 5160
rect 127066 5040 127072 5092
rect 127124 5080 127130 5092
rect 219710 5080 219716 5092
rect 127124 5052 219716 5080
rect 127124 5040 127130 5052
rect 219710 5040 219716 5052
rect 219768 5040 219774 5092
rect 248414 5040 248420 5092
rect 248472 5080 248478 5092
rect 501782 5080 501788 5092
rect 248472 5052 501788 5080
rect 248472 5040 248478 5052
rect 501782 5040 501788 5052
rect 501840 5040 501846 5092
rect 110506 4972 110512 5024
rect 110564 5012 110570 5024
rect 207934 5012 207940 5024
rect 110564 4984 207940 5012
rect 110564 4972 110570 4984
rect 207934 4972 207940 4984
rect 207992 4972 207998 5024
rect 251266 4972 251272 5024
rect 251324 5012 251330 5024
rect 537202 5012 537208 5024
rect 251324 4984 537208 5012
rect 251324 4972 251330 4984
rect 537202 4972 537208 4984
rect 537260 4972 537266 5024
rect 60826 4904 60832 4956
rect 60884 4944 60890 4956
rect 213914 4944 213920 4956
rect 60884 4916 213920 4944
rect 60884 4904 60890 4916
rect 213914 4904 213920 4916
rect 213972 4904 213978 4956
rect 230474 4904 230480 4956
rect 230532 4944 230538 4956
rect 239398 4944 239404 4956
rect 230532 4916 239404 4944
rect 230532 4904 230538 4916
rect 239398 4904 239404 4916
rect 239456 4904 239462 4956
rect 252646 4904 252652 4956
rect 252704 4944 252710 4956
rect 547874 4944 547880 4956
rect 252704 4916 547880 4944
rect 252704 4904 252710 4916
rect 547874 4904 547880 4916
rect 547932 4904 547938 4956
rect 15930 4836 15936 4888
rect 15988 4876 15994 4888
rect 42058 4876 42064 4888
rect 15988 4848 42064 4876
rect 15988 4836 15994 4848
rect 42058 4836 42064 4848
rect 42116 4836 42122 4888
rect 58434 4836 58440 4888
rect 58492 4876 58498 4888
rect 214006 4876 214012 4888
rect 58492 4848 214012 4876
rect 58492 4836 58498 4848
rect 214006 4836 214012 4848
rect 214064 4836 214070 4888
rect 214466 4836 214472 4888
rect 214524 4876 214530 4888
rect 226610 4876 226616 4888
rect 214524 4848 226616 4876
rect 214524 4836 214530 4848
rect 226610 4836 226616 4848
rect 226668 4836 226674 4888
rect 229554 4836 229560 4888
rect 229612 4876 229618 4888
rect 248782 4876 248788 4888
rect 229612 4848 248788 4876
rect 229612 4836 229618 4848
rect 248782 4836 248788 4848
rect 248840 4836 248846 4888
rect 252554 4836 252560 4888
rect 252612 4876 252618 4888
rect 551462 4876 551468 4888
rect 252612 4848 551468 4876
rect 252612 4836 252618 4848
rect 551462 4836 551468 4848
rect 551520 4836 551526 4888
rect 32398 4768 32404 4820
rect 32456 4808 32462 4820
rect 206278 4808 206284 4820
rect 32456 4780 206284 4808
rect 32456 4768 32462 4780
rect 206278 4768 206284 4780
rect 206336 4768 206342 4820
rect 210970 4768 210976 4820
rect 211028 4808 211034 4820
rect 226518 4808 226524 4820
rect 211028 4780 226524 4808
rect 211028 4768 211034 4780
rect 226518 4768 226524 4780
rect 226576 4768 226582 4820
rect 229646 4768 229652 4820
rect 229704 4808 229710 4820
rect 251174 4808 251180 4820
rect 229704 4780 251180 4808
rect 229704 4768 229710 4780
rect 251174 4768 251180 4780
rect 251232 4768 251238 4820
rect 255406 4768 255412 4820
rect 255464 4808 255470 4820
rect 578602 4808 578608 4820
rect 255464 4780 578608 4808
rect 255464 4768 255470 4780
rect 578602 4768 578608 4780
rect 578660 4768 578666 4820
rect 200298 4088 200304 4140
rect 200356 4128 200362 4140
rect 225690 4128 225696 4140
rect 200356 4100 225696 4128
rect 200356 4088 200362 4100
rect 225690 4088 225696 4100
rect 225748 4088 225754 4140
rect 185026 4020 185032 4072
rect 185084 4060 185090 4072
rect 210418 4060 210424 4072
rect 185084 4032 210424 4060
rect 185084 4020 185090 4032
rect 210418 4020 210424 4032
rect 210476 4020 210482 4072
rect 219250 4020 219256 4072
rect 219308 4060 219314 4072
rect 220814 4060 220820 4072
rect 219308 4032 220820 4060
rect 219308 4020 219314 4032
rect 220814 4020 220820 4032
rect 220872 4020 220878 4072
rect 177850 3952 177856 4004
rect 177908 3992 177914 4004
rect 204898 3992 204904 4004
rect 177908 3964 204904 3992
rect 177908 3952 177914 3964
rect 204898 3952 204904 3964
rect 204956 3952 204962 4004
rect 233878 3952 233884 4004
rect 233936 3992 233942 4004
rect 245194 3992 245200 4004
rect 233936 3964 245200 3992
rect 233936 3952 233942 3964
rect 245194 3952 245200 3964
rect 245252 3952 245258 4004
rect 132954 3884 132960 3936
rect 133012 3924 133018 3936
rect 187694 3924 187700 3936
rect 133012 3896 187700 3924
rect 133012 3884 133018 3896
rect 187694 3884 187700 3896
rect 187752 3884 187758 3936
rect 193214 3884 193220 3936
rect 193272 3924 193278 3936
rect 225046 3924 225052 3936
rect 193272 3896 225052 3924
rect 193272 3884 193278 3896
rect 225046 3884 225052 3896
rect 225104 3884 225110 3936
rect 229462 3884 229468 3936
rect 229520 3924 229526 3936
rect 242894 3924 242900 3936
rect 229520 3896 242900 3924
rect 229520 3884 229526 3896
rect 242894 3884 242900 3896
rect 242952 3884 242958 3936
rect 104526 3816 104532 3868
rect 104584 3856 104590 3868
rect 159358 3856 159364 3868
rect 104584 3828 159364 3856
rect 104584 3816 104590 3828
rect 159358 3816 159364 3828
rect 159416 3816 159422 3868
rect 166074 3816 166080 3868
rect 166132 3856 166138 3868
rect 201402 3856 201408 3868
rect 166132 3828 201408 3856
rect 166132 3816 166138 3828
rect 201402 3816 201408 3828
rect 201460 3816 201466 3868
rect 218054 3816 218060 3868
rect 218112 3856 218118 3868
rect 227346 3856 227352 3868
rect 218112 3828 227352 3856
rect 218112 3816 218118 3828
rect 227346 3816 227352 3828
rect 227404 3816 227410 3868
rect 229186 3816 229192 3868
rect 229244 3856 229250 3868
rect 239214 3856 239220 3868
rect 229244 3828 239220 3856
rect 229244 3816 229250 3828
rect 239214 3816 239220 3828
rect 239272 3816 239278 3868
rect 239398 3816 239404 3868
rect 239456 3856 239462 3868
rect 239456 3828 248414 3856
rect 239456 3816 239462 3828
rect 84470 3748 84476 3800
rect 84528 3788 84534 3800
rect 140038 3788 140044 3800
rect 84528 3760 140044 3788
rect 84528 3748 84534 3760
rect 140038 3748 140044 3760
rect 140096 3748 140102 3800
rect 168466 3748 168472 3800
rect 168524 3788 168530 3800
rect 213178 3788 213184 3800
rect 168524 3760 213184 3788
rect 168524 3748 168530 3760
rect 213178 3748 213184 3760
rect 213236 3748 213242 3800
rect 248386 3788 248414 3828
rect 257614 3816 257620 3868
rect 257672 3856 257678 3868
rect 264146 3856 264152 3868
rect 257672 3828 264152 3856
rect 257672 3816 257678 3828
rect 264146 3816 264152 3828
rect 264204 3816 264210 3868
rect 261754 3788 261760 3800
rect 248386 3760 261760 3788
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 276014 3748 276020 3800
rect 276072 3788 276078 3800
rect 276750 3788 276756 3800
rect 276072 3760 276756 3788
rect 276072 3748 276078 3760
rect 276750 3748 276756 3760
rect 276808 3748 276814 3800
rect 106918 3680 106924 3732
rect 106976 3720 106982 3732
rect 163498 3720 163504 3732
rect 106976 3692 163504 3720
rect 106976 3680 106982 3692
rect 163498 3680 163504 3692
rect 163556 3680 163562 3732
rect 179046 3680 179052 3732
rect 179104 3720 179110 3732
rect 224218 3720 224224 3732
rect 179104 3692 224224 3720
rect 179104 3680 179110 3692
rect 224218 3680 224224 3692
rect 224276 3680 224282 3732
rect 228266 3680 228272 3732
rect 228324 3720 228330 3732
rect 229830 3720 229836 3732
rect 228324 3692 229836 3720
rect 228324 3680 228330 3692
rect 229830 3680 229836 3692
rect 229888 3680 229894 3732
rect 296070 3720 296076 3732
rect 234586 3692 296076 3720
rect 99834 3612 99840 3664
rect 99892 3652 99898 3664
rect 156598 3652 156604 3664
rect 99892 3624 156604 3652
rect 99892 3612 99898 3624
rect 156598 3612 156604 3624
rect 156656 3612 156662 3664
rect 161290 3612 161296 3664
rect 161348 3652 161354 3664
rect 207658 3652 207664 3664
rect 161348 3624 207664 3652
rect 161348 3612 161354 3624
rect 207658 3612 207664 3624
rect 207716 3612 207722 3664
rect 216858 3612 216864 3664
rect 216916 3652 216922 3664
rect 222286 3652 222292 3664
rect 216916 3624 222292 3652
rect 216916 3612 216922 3624
rect 222286 3612 222292 3624
rect 222344 3612 222350 3664
rect 227898 3612 227904 3664
rect 227956 3652 227962 3664
rect 232222 3652 232228 3664
rect 227956 3624 232228 3652
rect 227956 3612 227962 3624
rect 232222 3612 232228 3624
rect 232280 3612 232286 3664
rect 233234 3612 233240 3664
rect 233292 3652 233298 3664
rect 234586 3652 234614 3692
rect 296070 3680 296076 3692
rect 296128 3680 296134 3732
rect 307846 3680 307852 3732
rect 307904 3720 307910 3732
rect 309042 3720 309048 3732
rect 307904 3692 309048 3720
rect 307904 3680 307910 3692
rect 309042 3680 309048 3692
rect 309100 3680 309106 3732
rect 316126 3680 316132 3732
rect 316184 3720 316190 3732
rect 317322 3720 317328 3732
rect 316184 3692 317328 3720
rect 316184 3680 316190 3692
rect 317322 3680 317328 3692
rect 317380 3680 317386 3732
rect 233292 3624 234614 3652
rect 233292 3612 233298 3624
rect 236638 3612 236644 3664
rect 236696 3652 236702 3664
rect 257062 3652 257068 3664
rect 236696 3624 257068 3652
rect 236696 3612 236702 3624
rect 257062 3612 257068 3624
rect 257120 3612 257126 3664
rect 257338 3612 257344 3664
rect 257396 3652 257402 3664
rect 458082 3652 458088 3664
rect 257396 3624 458088 3652
rect 257396 3612 257402 3624
rect 458082 3612 458088 3624
rect 458140 3612 458146 3664
rect 93854 3544 93860 3596
rect 93912 3584 93918 3596
rect 94774 3584 94780 3596
rect 93912 3556 94780 3584
rect 93912 3544 93918 3556
rect 94774 3544 94780 3556
rect 94832 3544 94838 3596
rect 102134 3544 102140 3596
rect 102192 3584 102198 3596
rect 103330 3584 103336 3596
rect 102192 3556 103336 3584
rect 102192 3544 102198 3556
rect 103330 3544 103336 3556
rect 103388 3544 103394 3596
rect 110414 3544 110420 3596
rect 110472 3584 110478 3596
rect 111610 3584 111616 3596
rect 110472 3556 111616 3584
rect 110472 3544 110478 3556
rect 111610 3544 111616 3556
rect 111668 3544 111674 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 209038 3584 209044 3596
rect 125928 3556 209044 3584
rect 125928 3544 125934 3556
rect 209038 3544 209044 3556
rect 209096 3544 209102 3596
rect 209774 3544 209780 3596
rect 209832 3584 209838 3596
rect 213270 3584 213276 3596
rect 209832 3556 213276 3584
rect 209832 3544 209838 3556
rect 213270 3544 213276 3556
rect 213328 3544 213334 3596
rect 229278 3544 229284 3596
rect 229336 3584 229342 3596
rect 253474 3584 253480 3596
rect 229336 3556 253480 3584
rect 229336 3544 229342 3556
rect 253474 3544 253480 3556
rect 253532 3544 253538 3596
rect 255958 3544 255964 3596
rect 256016 3584 256022 3596
rect 472250 3584 472256 3596
rect 256016 3556 472256 3584
rect 256016 3544 256022 3556
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 473354 3544 473360 3596
rect 473412 3584 473418 3596
rect 474182 3584 474188 3596
rect 473412 3556 474188 3584
rect 473412 3544 473418 3556
rect 474182 3544 474188 3556
rect 474240 3544 474246 3596
rect 484026 3584 484032 3596
rect 480226 3556 484032 3584
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20254 3516 20260 3528
rect 19392 3488 20260 3516
rect 19392 3476 19398 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 70302 3476 70308 3528
rect 70360 3516 70366 3528
rect 70360 3488 125364 3516
rect 70360 3476 70366 3488
rect 30098 3408 30104 3460
rect 30156 3448 30162 3460
rect 125336 3448 125364 3488
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128170 3516 128176 3528
rect 127032 3488 128176 3516
rect 127032 3476 127038 3488
rect 128170 3476 128176 3488
rect 128228 3476 128234 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 219526 3516 219532 3528
rect 129424 3488 219532 3516
rect 129424 3476 129430 3488
rect 219526 3476 219532 3488
rect 219584 3476 219590 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 228174 3516 228180 3528
rect 226392 3488 228180 3516
rect 226392 3476 226398 3488
rect 228174 3476 228180 3488
rect 228232 3476 228238 3528
rect 230106 3476 230112 3528
rect 230164 3516 230170 3528
rect 244090 3516 244096 3528
rect 230164 3488 244096 3516
rect 230164 3476 230170 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 248046 3476 248052 3528
rect 248104 3516 248110 3528
rect 480226 3516 480254 3556
rect 484026 3544 484032 3556
rect 484084 3544 484090 3596
rect 248104 3488 480254 3516
rect 248104 3476 248110 3488
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 127618 3448 127624 3460
rect 30156 3420 122834 3448
rect 125336 3420 127624 3448
rect 30156 3408 30162 3420
rect 122806 3312 122834 3420
rect 127618 3408 127624 3420
rect 127676 3408 127682 3460
rect 207750 3448 207756 3460
rect 132466 3420 207756 3448
rect 132466 3312 132494 3420
rect 207750 3408 207756 3420
rect 207808 3408 207814 3460
rect 229370 3408 229376 3460
rect 229428 3448 229434 3460
rect 246390 3448 246396 3460
rect 229428 3420 246396 3448
rect 229428 3408 229434 3420
rect 246390 3408 246396 3420
rect 246448 3408 246454 3460
rect 252462 3408 252468 3460
rect 252520 3448 252526 3460
rect 530118 3448 530124 3460
rect 252520 3420 530124 3448
rect 252520 3408 252526 3420
rect 530118 3408 530124 3420
rect 530176 3408 530182 3460
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169570 3380 169576 3392
rect 168432 3352 169576 3380
rect 168432 3340 168438 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186130 3380 186136 3392
rect 184992 3352 186136 3380
rect 184992 3340 184998 3352
rect 186130 3340 186136 3352
rect 186188 3340 186194 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 207842 3380 207848 3392
rect 190880 3352 207848 3380
rect 190880 3340 190886 3352
rect 207842 3340 207848 3352
rect 207900 3340 207906 3392
rect 227990 3340 227996 3392
rect 228048 3380 228054 3392
rect 231026 3380 231032 3392
rect 228048 3352 231032 3380
rect 228048 3340 228054 3352
rect 231026 3340 231032 3352
rect 231084 3340 231090 3392
rect 231118 3340 231124 3392
rect 231176 3380 231182 3392
rect 237006 3380 237012 3392
rect 231176 3352 237012 3380
rect 231176 3340 231182 3352
rect 237006 3340 237012 3352
rect 237064 3340 237070 3392
rect 239214 3340 239220 3392
rect 239272 3380 239278 3392
rect 247586 3380 247592 3392
rect 239272 3352 247592 3380
rect 239272 3340 239278 3352
rect 247586 3340 247592 3352
rect 247644 3340 247650 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365806 3340 365812 3392
rect 365864 3380 365870 3392
rect 367002 3380 367008 3392
rect 365864 3352 367008 3380
rect 365864 3340 365870 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 122806 3284 132494 3312
rect 223942 3136 223948 3188
rect 224000 3176 224006 3188
rect 228082 3176 228088 3188
rect 224000 3148 228088 3176
rect 224000 3136 224006 3148
rect 228082 3136 228088 3148
rect 228140 3136 228146 3188
rect 213362 3000 213368 3052
rect 213420 3040 213426 3052
rect 220078 3040 220084 3052
rect 213420 3012 220084 3040
rect 213420 3000 213426 3012
rect 220078 3000 220084 3012
rect 220136 3000 220142 3052
rect 221550 3000 221556 3052
rect 221608 3040 221614 3052
rect 227162 3040 227168 3052
rect 221608 3012 227168 3040
rect 221608 3000 221614 3012
rect 227162 3000 227168 3012
rect 227220 3000 227226 3052
rect 249978 3000 249984 3052
rect 250036 3040 250042 3052
rect 256694 3040 256700 3052
rect 250036 3012 256700 3040
rect 250036 3000 250042 3012
rect 256694 3000 256700 3012
rect 256752 3000 256758 3052
rect 225138 2932 225144 2984
rect 225196 2972 225202 2984
rect 226426 2972 226432 2984
rect 225196 2944 226432 2972
rect 225196 2932 225202 2944
rect 226426 2932 226432 2944
rect 226484 2932 226490 2984
rect 423674 1640 423680 1692
rect 423732 1680 423738 1692
rect 424962 1680 424968 1692
rect 423732 1652 424968 1680
rect 423732 1640 423738 1652
rect 424962 1640 424968 1652
rect 425020 1640 425026 1692
rect 448514 1640 448520 1692
rect 448572 1680 448578 1692
rect 449802 1680 449808 1692
rect 448572 1652 449808 1680
rect 448572 1640 448578 1652
rect 449802 1640 449808 1652
rect 449860 1640 449866 1692
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 154120 700476 154172 700528
rect 177396 700476 177448 700528
rect 402244 700476 402296 700528
rect 429844 700476 429896 700528
rect 137836 700408 137888 700460
rect 173256 700408 173308 700460
rect 188988 700408 189040 700460
rect 202788 700408 202840 700460
rect 298836 700408 298888 700460
rect 332508 700408 332560 700460
rect 402336 700408 402388 700460
rect 462320 700408 462372 700460
rect 24308 700340 24360 700392
rect 33784 700340 33836 700392
rect 40500 700340 40552 700392
rect 51724 700340 51776 700392
rect 105452 700340 105504 700392
rect 177304 700340 177356 700392
rect 190000 700340 190052 700392
rect 218980 700340 219032 700392
rect 290556 700340 290608 700392
rect 348792 700340 348844 700392
rect 392584 700340 392636 700392
rect 478512 700340 478564 700392
rect 8116 700272 8168 700324
rect 55864 700272 55916 700324
rect 89168 700272 89220 700324
rect 171784 700272 171836 700324
rect 189908 700272 189960 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 281540 700272 281592 700324
rect 294604 700272 294656 700324
rect 364984 700272 365036 700324
rect 393964 700272 394016 700324
rect 494796 700272 494848 700324
rect 505744 700272 505796 700324
rect 559656 700272 559708 700324
rect 170312 699660 170364 699712
rect 173164 699660 173216 699712
rect 298744 699660 298796 699712
rect 300124 699660 300176 699712
rect 409144 699660 409196 699712
rect 413652 699660 413704 699712
rect 290464 696940 290516 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 15844 683136 15896 683188
rect 533344 683136 533396 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 37924 670692 37976 670744
rect 502984 670692 503036 670744
rect 580172 670692 580224 670744
rect 2780 656956 2832 657008
rect 4804 656956 4856 657008
rect 503076 643084 503128 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 51816 632068 51868 632120
rect 523684 630640 523736 630692
rect 580172 630640 580224 630692
rect 503168 616836 503220 616888
rect 580172 616836 580224 616888
rect 3148 605888 3200 605940
rect 6184 605888 6236 605940
rect 407764 600244 407816 600296
rect 407948 600244 408000 600296
rect 78128 599972 78180 600024
rect 187240 599972 187292 600024
rect 297824 599972 297876 600024
rect 408224 599972 408276 600024
rect 78036 599904 78088 599956
rect 187148 599904 187200 599956
rect 78220 599836 78272 599888
rect 187332 599836 187384 599888
rect 78588 599768 78640 599820
rect 186596 599768 186648 599820
rect 297364 599768 297416 599820
rect 297824 599768 297876 599820
rect 78404 599700 78456 599752
rect 187056 599700 187108 599752
rect 78496 599632 78548 599684
rect 186872 599632 186924 599684
rect 297916 599564 297968 599616
rect 407764 599564 407816 599616
rect 297272 599360 297324 599412
rect 297916 599360 297968 599412
rect 297456 598884 297508 598936
rect 407580 598884 407632 598936
rect 297548 598816 297600 598868
rect 407396 598816 407448 598868
rect 297180 598272 297232 598324
rect 298008 598272 298060 598324
rect 407488 598204 407540 598256
rect 115848 597524 115900 597576
rect 225512 597524 225564 597576
rect 282368 597524 282420 597576
rect 335360 597524 335412 597576
rect 444380 597524 444432 597576
rect 126888 597456 126940 597508
rect 234620 597456 234672 597508
rect 326160 597456 326212 597508
rect 434720 597456 434772 597508
rect 136548 597388 136600 597440
rect 245476 597388 245528 597440
rect 111708 597320 111760 597372
rect 219440 597320 219492 597372
rect 220728 597320 220780 597372
rect 103152 597252 103204 597304
rect 212356 597252 212408 597304
rect 140688 597184 140740 597236
rect 131028 597116 131080 597168
rect 106188 597048 106240 597100
rect 215300 597048 215352 597100
rect 121368 596980 121420 597032
rect 100668 596912 100720 596964
rect 209964 596912 210016 596964
rect 211068 596912 211120 596964
rect 103428 596844 103480 596896
rect 213828 596844 213880 596896
rect 104808 596776 104860 596828
rect 214840 596776 214892 596828
rect 281632 597388 281684 597440
rect 350448 597388 350500 597440
rect 459560 597388 459612 597440
rect 330392 597320 330444 597372
rect 440240 597320 440292 597372
rect 281724 597252 281776 597304
rect 345664 597252 345716 597304
rect 455420 597252 455472 597304
rect 282184 597184 282236 597236
rect 340512 597184 340564 597236
rect 449900 597184 449952 597236
rect 282092 597116 282144 597168
rect 250536 597048 250588 597100
rect 284300 597048 284352 597100
rect 323400 597116 323452 597168
rect 433340 597116 433392 597168
rect 324320 597048 324372 597100
rect 324780 597048 324832 597100
rect 434720 597048 434772 597100
rect 281908 596980 281960 597032
rect 360568 596980 360620 597032
rect 240508 596912 240560 596964
rect 281632 596912 281684 596964
rect 282000 596912 282052 596964
rect 284668 596912 284720 596964
rect 299388 596912 299440 596964
rect 314660 596912 314712 596964
rect 470600 596912 470652 596964
rect 234620 596844 234672 596896
rect 281724 596844 281776 596896
rect 282276 596844 282328 596896
rect 319996 596844 320048 596896
rect 429200 596844 429252 596896
rect 230664 596776 230716 596828
rect 282184 596776 282236 596828
rect 284944 596776 284996 596828
rect 322296 596776 322348 596828
rect 431960 596776 432012 596828
rect 220728 596708 220780 596760
rect 280988 596708 281040 596760
rect 330392 596708 330444 596760
rect 354680 596708 354732 596760
rect 465080 596708 465132 596760
rect 215300 596640 215352 596692
rect 284576 596640 284628 596692
rect 214840 596572 214892 596624
rect 284484 596572 284536 596624
rect 324320 596572 324372 596624
rect 213828 596504 213880 596556
rect 284300 596504 284352 596556
rect 284576 596504 284628 596556
rect 326160 596504 326212 596556
rect 212448 596436 212500 596488
rect 284392 596436 284444 596488
rect 211068 596368 211120 596420
rect 282276 596368 282328 596420
rect 79784 596300 79836 596352
rect 92480 596300 92532 596352
rect 188712 596300 188764 596352
rect 202880 596300 202932 596352
rect 209044 596300 209096 596352
rect 282000 596300 282052 596352
rect 282092 596300 282144 596352
rect 408224 596300 408276 596352
rect 422576 596300 422628 596352
rect 79876 596232 79928 596284
rect 94044 596232 94096 596284
rect 188896 596232 188948 596284
rect 204352 596232 204404 596284
rect 207664 596232 207716 596284
rect 284760 596232 284812 596284
rect 299296 596232 299348 596284
rect 311900 596232 311952 596284
rect 407948 596232 408000 596284
rect 423680 596232 423732 596284
rect 79968 596164 80020 596216
rect 95240 596164 95292 596216
rect 188804 596164 188856 596216
rect 204260 596164 204312 596216
rect 212356 596164 212408 596216
rect 284944 596164 284996 596216
rect 299204 596164 299256 596216
rect 313280 596164 313332 596216
rect 407764 596164 407816 596216
rect 425060 596164 425112 596216
rect 281632 591336 281684 591388
rect 282000 591336 282052 591388
rect 281632 591200 281684 591252
rect 282368 591200 282420 591252
rect 283564 590656 283616 590708
rect 579804 590656 579856 590708
rect 78312 584400 78364 584452
rect 186688 584400 186740 584452
rect 2780 579912 2832 579964
rect 4896 579912 4948 579964
rect 501604 563048 501656 563100
rect 580172 563048 580224 563100
rect 3332 553528 3384 553580
rect 7564 553528 7616 553580
rect 515404 536800 515456 536852
rect 579896 536800 579948 536852
rect 2780 527212 2832 527264
rect 4988 527212 5040 527264
rect 284944 526396 284996 526448
rect 297180 526396 297232 526448
rect 297732 526396 297784 526448
rect 294696 525920 294748 525972
rect 297272 525920 297324 525972
rect 298008 525920 298060 525972
rect 186872 525852 186924 525904
rect 187700 525852 187752 525904
rect 519544 524424 519596 524476
rect 580172 524424 580224 524476
rect 285588 523744 285640 523796
rect 297364 523744 297416 523796
rect 298008 523744 298060 523796
rect 284208 523676 284260 523728
rect 297640 523676 297692 523728
rect 297916 523676 297968 523728
rect 187516 521568 187568 521620
rect 188160 521568 188212 521620
rect 284116 520956 284168 521008
rect 297456 520956 297508 521008
rect 284024 520888 284076 520940
rect 297824 520888 297876 520940
rect 187148 518372 187200 518424
rect 188068 518372 188120 518424
rect 282828 518168 282880 518220
rect 297548 518168 297600 518220
rect 3332 514768 3384 514820
rect 14464 514768 14516 514820
rect 549904 510620 549956 510672
rect 580172 510620 580224 510672
rect 3332 500964 3384 501016
rect 15936 500964 15988 501016
rect 78128 489812 78180 489864
rect 187976 489812 188028 489864
rect 408132 489812 408184 489864
rect 78036 489744 78088 489796
rect 188068 489744 188120 489796
rect 284024 489744 284076 489796
rect 284208 489744 284260 489796
rect 407672 489744 407724 489796
rect 77760 489676 77812 489728
rect 188160 489676 188212 489728
rect 284116 489676 284168 489728
rect 407580 489676 407632 489728
rect 78312 489608 78364 489660
rect 188344 489608 188396 489660
rect 297916 489608 297968 489660
rect 408408 489608 408460 489660
rect 77576 489540 77628 489592
rect 187792 489540 187844 489592
rect 297824 489540 297876 489592
rect 407856 489540 407908 489592
rect 78496 489472 78548 489524
rect 187700 489472 187752 489524
rect 77668 489404 77720 489456
rect 187056 489404 187108 489456
rect 78588 489336 78640 489388
rect 186964 489336 187016 489388
rect 188344 489132 188396 489184
rect 240784 489132 240836 489184
rect 187976 488860 188028 488912
rect 188620 488860 188672 488912
rect 110512 488792 110564 488844
rect 220728 488792 220780 488844
rect 187792 488724 187844 488776
rect 188252 488724 188304 488776
rect 215300 488724 215352 488776
rect 242900 488724 242952 488776
rect 325332 488724 325384 488776
rect 120632 488656 120684 488708
rect 230480 488656 230532 488708
rect 231768 488656 231820 488708
rect 283656 488656 283708 488708
rect 284208 488656 284260 488708
rect 297364 488656 297416 488708
rect 297824 488656 297876 488708
rect 336648 488724 336700 488776
rect 444380 488724 444432 488776
rect 434720 488656 434772 488708
rect 115664 488588 115716 488640
rect 226248 488588 226300 488640
rect 335452 488588 335504 488640
rect 336648 488588 336700 488640
rect 340604 488588 340656 488640
rect 449900 488588 449952 488640
rect 105360 488520 105412 488572
rect 215300 488520 215352 488572
rect 220728 488520 220780 488572
rect 330484 488520 330536 488572
rect 440240 488520 440292 488572
rect 79784 488452 79836 488504
rect 92940 488452 92992 488504
rect 188712 488452 188764 488504
rect 231768 488452 231820 488504
rect 340604 488452 340656 488504
rect 407948 488452 408000 488504
rect 423680 488452 423732 488504
rect 79876 488384 79928 488436
rect 94228 488384 94280 488436
rect 188804 488384 188856 488436
rect 408224 488384 408276 488436
rect 422576 488384 422628 488436
rect 79968 488316 80020 488368
rect 95332 488316 95384 488368
rect 312544 488180 312596 488232
rect 408224 488180 408276 488232
rect 318892 488112 318944 488164
rect 427820 488112 427872 488164
rect 188712 488044 188764 488096
rect 202880 488044 202932 488096
rect 326344 488044 326396 488096
rect 434720 488044 434772 488096
rect 188804 487976 188856 488028
rect 204260 487976 204312 488028
rect 360476 487976 360528 488028
rect 470600 487976 470652 488028
rect 102416 487908 102468 487960
rect 211804 487908 211856 487960
rect 219624 487908 219676 487960
rect 281540 487908 281592 487960
rect 345756 487908 345808 487960
rect 455420 487908 455472 487960
rect 135536 487840 135588 487892
rect 244556 487840 244608 487892
rect 355784 487840 355836 487892
rect 465080 487840 465132 487892
rect 125600 487772 125652 487824
rect 235632 487772 235684 487824
rect 235908 487772 235960 487824
rect 97816 487704 97868 487756
rect 207664 487704 207716 487756
rect 105728 487636 105780 487688
rect 215944 487636 215996 487688
rect 104808 487568 104860 487620
rect 214564 487568 214616 487620
rect 99196 487500 99248 487552
rect 209044 487500 209096 487552
rect 100024 487432 100076 487484
rect 210056 487432 210108 487484
rect 211068 487432 211120 487484
rect 241428 487772 241480 487824
rect 350356 487772 350408 487824
rect 459560 487772 459612 487824
rect 318064 487704 318116 487756
rect 426440 487704 426492 487756
rect 320824 487636 320876 487688
rect 430580 487636 430632 487688
rect 320088 487568 320140 487620
rect 429200 487568 429252 487620
rect 322204 487500 322256 487552
rect 432052 487500 432104 487552
rect 345756 487432 345808 487484
rect 103428 487364 103480 487416
rect 213184 487364 213236 487416
rect 101128 487296 101180 487348
rect 211160 487296 211212 487348
rect 212448 487296 212500 487348
rect 140688 487228 140740 487280
rect 250444 487364 250496 487416
rect 251088 487364 251140 487416
rect 360476 487364 360528 487416
rect 244556 487296 244608 487348
rect 245568 487296 245620 487348
rect 355784 487296 355836 487348
rect 323584 487228 323636 487280
rect 433340 487228 433392 487280
rect 130660 487160 130712 487212
rect 241428 487160 241480 487212
rect 324320 487160 324372 487212
rect 324872 487160 324924 487212
rect 434720 487160 434772 487212
rect 212448 486480 212500 486532
rect 247684 486480 247736 486532
rect 187700 486412 187752 486464
rect 241520 486412 241572 486464
rect 244924 486412 244976 486464
rect 318892 486412 318944 486464
rect 187056 485052 187108 485104
rect 261484 485052 261536 485104
rect 261576 485052 261628 485104
rect 297916 485052 297968 485104
rect 211160 484372 211212 484424
rect 580172 484372 580224 484424
rect 241520 484304 241572 484356
rect 284944 484304 284996 484356
rect 242808 482332 242860 482384
rect 294696 482332 294748 482384
rect 211068 482264 211120 482316
rect 246120 482264 246172 482316
rect 250352 482264 250404 482316
rect 324320 482264 324372 482316
rect 207664 481040 207716 481092
rect 243544 481040 243596 481092
rect 240140 480972 240192 481024
rect 284116 480972 284168 481024
rect 236000 480904 236052 480956
rect 297456 480904 297508 480956
rect 239956 479544 240008 479596
rect 284024 479544 284076 479596
rect 220728 479476 220780 479528
rect 244280 479476 244332 479528
rect 251640 479476 251692 479528
rect 326344 479476 326396 479528
rect 189080 478796 189132 478848
rect 241888 478796 241940 478848
rect 245844 478796 245896 478848
rect 319444 478796 319496 478848
rect 240048 478184 240100 478236
rect 282368 478184 282420 478236
rect 188252 478116 188304 478168
rect 240876 478116 240928 478168
rect 241888 477980 241940 478032
rect 242808 477980 242860 478032
rect 188620 477436 188672 477488
rect 240140 477436 240192 477488
rect 245568 477436 245620 477488
rect 249800 477436 249852 477488
rect 187608 476756 187660 476808
rect 236368 476756 236420 476808
rect 249156 476756 249208 476808
rect 323584 476756 323636 476808
rect 299112 476416 299164 476468
rect 299388 476416 299440 476468
rect 214564 476008 214616 476060
rect 250352 476008 250404 476060
rect 298652 476008 298704 476060
rect 299204 476008 299256 476060
rect 313924 476008 313976 476060
rect 173256 475464 173308 475516
rect 221096 475464 221148 475516
rect 51816 475396 51868 475448
rect 224132 475396 224184 475448
rect 238116 475396 238168 475448
rect 298652 475396 298704 475448
rect 15844 475328 15896 475380
rect 224040 475328 224092 475380
rect 249064 475328 249116 475380
rect 322204 475328 322256 475380
rect 3056 474716 3108 474768
rect 14556 474716 14608 474768
rect 188528 474648 188580 474700
rect 238760 474648 238812 474700
rect 239956 474648 240008 474700
rect 247040 474648 247092 474700
rect 247684 474648 247736 474700
rect 320824 474648 320876 474700
rect 299388 474580 299440 474632
rect 312544 474580 312596 474632
rect 238024 473968 238076 474020
rect 299388 473968 299440 474020
rect 188344 473288 188396 473340
rect 239128 473288 239180 473340
rect 240048 473288 240100 473340
rect 243084 473288 243136 473340
rect 243544 473288 243596 473340
rect 318064 473288 318116 473340
rect 241428 472676 241480 472728
rect 248696 472676 248748 472728
rect 218060 472608 218112 472660
rect 290556 472608 290608 472660
rect 215944 471928 215996 471980
rect 251640 471928 251692 471980
rect 298652 471928 298704 471980
rect 299112 471928 299164 471980
rect 315304 471928 315356 471980
rect 177396 471248 177448 471300
rect 221280 471248 221332 471300
rect 238208 471248 238260 471300
rect 298652 471248 298704 471300
rect 217324 470568 217376 470620
rect 580172 470568 580224 470620
rect 216864 469888 216916 469940
rect 392584 469888 392636 469940
rect 216680 469820 216732 469872
rect 402336 469820 402388 469872
rect 186964 469140 187016 469192
rect 261208 469140 261260 469192
rect 261208 468868 261260 468920
rect 261576 468868 261628 468920
rect 213920 468528 213972 468580
rect 523684 468528 523736 468580
rect 215300 468460 215352 468512
rect 533344 468460 533396 468512
rect 218244 467236 218296 467288
rect 298836 467236 298888 467288
rect 77944 467168 77996 467220
rect 236184 467168 236236 467220
rect 214104 467100 214156 467152
rect 580264 467100 580316 467152
rect 218152 465740 218204 465792
rect 397460 465740 397512 465792
rect 215484 465672 215536 465724
rect 527180 465672 527232 465724
rect 218336 464448 218388 464500
rect 409144 464448 409196 464500
rect 214196 464380 214248 464432
rect 503076 464380 503128 464432
rect 212540 464312 212592 464364
rect 515404 464312 515456 464364
rect 51724 463088 51776 463140
rect 222660 463088 222712 463140
rect 236276 463088 236328 463140
rect 408040 463088 408092 463140
rect 216956 463020 217008 463072
rect 402244 463020 402296 463072
rect 212724 462952 212776 463004
rect 549904 462952 549956 463004
rect 3424 462340 3476 462392
rect 226984 462340 227036 462392
rect 217048 461796 217100 461848
rect 393964 461796 394016 461848
rect 3516 461728 3568 461780
rect 225604 461728 225656 461780
rect 215576 461660 215628 461712
rect 505744 461660 505796 461712
rect 216772 461592 216824 461644
rect 542360 461592 542412 461644
rect 215392 460300 215444 460352
rect 502984 460300 503036 460352
rect 214380 460232 214432 460284
rect 503168 460232 503220 460284
rect 212816 460164 212868 460216
rect 519544 460164 519596 460216
rect 213184 459484 213236 459536
rect 248972 459484 249024 459536
rect 249156 459484 249208 459536
rect 204904 459416 204956 459468
rect 238208 459416 238260 459468
rect 205088 459348 205140 459400
rect 238116 459348 238168 459400
rect 237932 458872 237984 458924
rect 238208 458872 238260 458924
rect 246304 458872 246356 458924
rect 371516 458872 371568 458924
rect 260932 458804 260984 458856
rect 309048 458804 309100 458856
rect 298836 458736 298888 458788
rect 329656 458736 329708 458788
rect 295984 458668 296036 458720
rect 346400 458668 346452 458720
rect 298928 458600 298980 458652
rect 354772 458600 354824 458652
rect 299572 458532 299624 458584
rect 359280 458532 359332 458584
rect 260196 458464 260248 458516
rect 321284 458464 321336 458516
rect 297548 458396 297600 458448
rect 363144 458396 363196 458448
rect 299020 458328 299072 458380
rect 367652 458328 367704 458380
rect 237840 458260 237892 458312
rect 238116 458260 238168 458312
rect 254584 458260 254636 458312
rect 379888 458260 379940 458312
rect 14464 457580 14516 457632
rect 227076 457580 227128 457632
rect 3608 457512 3660 457564
rect 224960 457512 225012 457564
rect 213552 457444 213604 457496
rect 501604 457444 501656 457496
rect 241796 457240 241848 457292
rect 312912 457240 312964 457292
rect 232136 457172 232188 457224
rect 325792 457172 325844 457224
rect 243636 457104 243688 457156
rect 338028 457104 338080 457156
rect 242992 457036 243044 457088
rect 342536 457036 342588 457088
rect 232596 456968 232648 457020
rect 334164 456968 334216 457020
rect 241704 456900 241756 456952
rect 350908 456900 350960 456952
rect 231124 456832 231176 456884
rect 376024 456832 376076 456884
rect 211344 456764 211396 456816
rect 580172 456764 580224 456816
rect 223212 456220 223264 456272
rect 317420 456220 317472 456272
rect 258080 456152 258132 456204
rect 385316 456152 385368 456204
rect 255780 456084 255832 456136
rect 384120 456084 384172 456136
rect 250076 456016 250128 456068
rect 384212 456016 384264 456068
rect 244740 455948 244792 456000
rect 384028 455948 384080 456000
rect 239036 455880 239088 455932
rect 385040 455880 385092 455932
rect 238944 455812 238996 455864
rect 385408 455812 385460 455864
rect 237564 455744 237616 455796
rect 385224 455744 385276 455796
rect 224960 455676 225012 455728
rect 225420 455676 225472 455728
rect 385500 455676 385552 455728
rect 299664 455608 299716 455660
rect 385132 455608 385184 455660
rect 211528 455540 211580 455592
rect 384304 455540 384356 455592
rect 224040 455472 224092 455524
rect 383568 455472 383620 455524
rect 211436 455404 211488 455456
rect 580264 455404 580316 455456
rect 37924 455336 37976 455388
rect 223764 455336 223816 455388
rect 224040 455336 224092 455388
rect 299848 455336 299900 455388
rect 304172 455336 304224 455388
rect 215668 454792 215720 454844
rect 290464 454792 290516 454844
rect 15936 454724 15988 454776
rect 226616 454724 226668 454776
rect 254492 454724 254544 454776
rect 299848 454724 299900 454776
rect 7564 454656 7616 454708
rect 225512 454656 225564 454708
rect 252560 454656 252612 454708
rect 299572 454656 299624 454708
rect 214012 453500 214064 453552
rect 283564 453500 283616 453552
rect 219532 453432 219584 453484
rect 298744 453432 298796 453484
rect 71780 453364 71832 453416
rect 222292 453364 222344 453416
rect 4804 453296 4856 453348
rect 223580 453296 223632 453348
rect 248604 453296 248656 453348
rect 297548 453296 297600 453348
rect 240784 452548 240836 452600
rect 285036 452548 285088 452600
rect 177304 452072 177356 452124
rect 221004 452072 221056 452124
rect 55864 452004 55916 452056
rect 222384 452004 222436 452056
rect 14556 451936 14608 451988
rect 226892 451936 226944 451988
rect 4988 451868 5040 451920
rect 225144 451868 225196 451920
rect 226248 451868 226300 451920
rect 245752 451868 245804 451920
rect 248052 451868 248104 451920
rect 299756 451868 299808 451920
rect 240324 451256 240376 451308
rect 298008 451256 298060 451308
rect 240876 451188 240928 451240
rect 283656 451188 283708 451240
rect 241704 451052 241756 451104
rect 241980 451052 242032 451104
rect 173164 450712 173216 450764
rect 221096 450712 221148 450764
rect 218704 450644 218756 450696
rect 294604 450644 294656 450696
rect 6184 450576 6236 450628
rect 224776 450576 224828 450628
rect 4896 450508 4948 450560
rect 225328 450508 225380 450560
rect 259828 450508 259880 450560
rect 299020 450508 299072 450560
rect 240692 449896 240744 449948
rect 240876 449896 240928 449948
rect 211804 449828 211856 449880
rect 248512 449828 248564 449880
rect 259552 449828 259604 449880
rect 284484 449828 284536 449880
rect 209044 449760 209096 449812
rect 245016 449760 245068 449812
rect 257896 449760 257948 449812
rect 282000 449760 282052 449812
rect 258632 449692 258684 449744
rect 284300 449692 284352 449744
rect 255688 449624 255740 449676
rect 282184 449624 282236 449676
rect 257344 449556 257396 449608
rect 284852 449556 284904 449608
rect 255136 449488 255188 449540
rect 282276 449488 282328 449540
rect 248512 449420 248564 449472
rect 249064 449420 249116 449472
rect 253480 449420 253532 449472
rect 280988 449420 281040 449472
rect 256240 449352 256292 449404
rect 284392 449352 284444 449404
rect 252376 449284 252428 449336
rect 281816 449284 281868 449336
rect 254308 449216 254360 449268
rect 298928 449216 298980 449268
rect 253756 449148 253808 449200
rect 298836 449148 298888 449200
rect 260656 449080 260708 449132
rect 284576 449080 284628 449132
rect 259000 449012 259052 449064
rect 282092 449012 282144 449064
rect 260104 448944 260156 448996
rect 281908 448944 281960 448996
rect 33784 448468 33836 448520
rect 223212 448468 223264 448520
rect 261484 448468 261536 448520
rect 267096 448468 267148 448520
rect 297364 448468 297416 448520
rect 203524 448400 203576 448452
rect 237472 448400 237524 448452
rect 238024 448400 238076 448452
rect 171784 447856 171836 447908
rect 222568 447856 222620 447908
rect 235908 447856 235960 447908
rect 247960 447856 248012 447908
rect 2872 447788 2924 447840
rect 227260 447788 227312 447840
rect 231768 447788 231820 447840
rect 246856 447788 246908 447840
rect 252100 447788 252152 447840
rect 295984 447788 296036 447840
rect 218060 447312 218112 447364
rect 219072 447312 219124 447364
rect 225420 447312 225472 447364
rect 225696 447312 225748 447364
rect 236000 447312 236052 447364
rect 236460 447312 236512 447364
rect 218244 447244 218296 447296
rect 218796 447244 218848 447296
rect 221004 447244 221056 447296
rect 221832 447244 221884 447296
rect 225144 447244 225196 447296
rect 225972 447244 226024 447296
rect 236276 447244 236328 447296
rect 236736 447244 236788 447296
rect 247684 447108 247736 447160
rect 297364 447108 297416 447160
rect 226708 446836 226760 446888
rect 227076 446836 227128 446888
rect 265900 446836 265952 446888
rect 212632 446768 212684 446820
rect 217324 446768 217376 446820
rect 225052 446768 225104 446820
rect 225604 446768 225656 446820
rect 264704 446768 264756 446820
rect 211160 446700 211212 446752
rect 212356 446700 212408 446752
rect 212540 446700 212592 446752
rect 213184 446700 213236 446752
rect 229468 446700 229520 446752
rect 264520 446700 264572 446752
rect 204904 446632 204956 446684
rect 231400 446632 231452 446684
rect 247132 446632 247184 446684
rect 299204 446632 299256 446684
rect 211436 446564 211488 446616
rect 211804 446564 211856 446616
rect 212816 446564 212868 446616
rect 213460 446564 213512 446616
rect 213920 446564 213972 446616
rect 215116 446564 215168 446616
rect 215576 446564 215628 446616
rect 216220 446564 216272 446616
rect 216680 446564 216732 446616
rect 217324 446564 217376 446616
rect 229008 446564 229060 446616
rect 251732 446564 251784 446616
rect 256792 446564 256844 446616
rect 281724 446564 281776 446616
rect 6184 446496 6236 446548
rect 230848 446496 230900 446548
rect 237932 446496 237984 446548
rect 238576 446496 238628 446548
rect 238944 446496 238996 446548
rect 239956 446496 240008 446548
rect 241520 446496 241572 446548
rect 242440 446496 242492 446548
rect 244372 446496 244424 446548
rect 246304 446496 246356 446548
rect 254400 446496 254452 446548
rect 281632 446496 281684 446548
rect 188988 446428 189040 446480
rect 220636 446428 220688 446480
rect 229100 446428 229152 446480
rect 260840 446428 260892 446480
rect 190000 446360 190052 446412
rect 220912 446360 220964 446412
rect 222568 446360 222620 446412
rect 229652 446360 229704 446412
rect 229744 446360 229796 446412
rect 258448 446360 258500 446412
rect 261760 446360 261812 446412
rect 299848 446360 299900 446412
rect 200856 446292 200908 446344
rect 228364 446292 228416 446344
rect 242900 446292 242952 446344
rect 243544 446292 243596 446344
rect 202420 446224 202472 446276
rect 233056 446224 233108 446276
rect 241612 446224 241664 446276
rect 257436 446224 257488 446276
rect 184204 446156 184256 446208
rect 229192 446156 229244 446208
rect 206560 446088 206612 446140
rect 247500 446088 247552 446140
rect 257620 446088 257672 446140
rect 299388 446088 299440 446140
rect 208216 446020 208268 446072
rect 251824 446020 251876 446072
rect 255412 446020 255464 446072
rect 298652 446020 298704 446072
rect 211252 445952 211304 446004
rect 299296 445952 299348 446004
rect 209872 445884 209924 445936
rect 299020 445884 299072 445936
rect 14464 445816 14516 445868
rect 230020 445816 230072 445868
rect 253204 445816 253256 445868
rect 297364 445816 297416 445868
rect 204168 445748 204220 445800
rect 232228 445748 232280 445800
rect 249892 445748 249944 445800
rect 254584 445748 254636 445800
rect 250076 445544 250128 445596
rect 250996 445544 251048 445596
rect 6276 445408 6328 445460
rect 229468 445408 229520 445460
rect 238760 445408 238812 445460
rect 239680 445408 239732 445460
rect 243084 445408 243136 445460
rect 244096 445408 244148 445460
rect 106924 445340 106976 445392
rect 228548 445340 228600 445392
rect 248972 445340 249024 445392
rect 249616 445340 249668 445392
rect 203616 445272 203668 445324
rect 231124 445272 231176 445324
rect 237564 445272 237616 445324
rect 238300 445272 238352 445324
rect 202328 445204 202380 445256
rect 233608 445204 233660 445256
rect 241796 445204 241848 445256
rect 242716 445204 242768 445256
rect 200764 445136 200816 445188
rect 232596 445136 232648 445188
rect 232780 445136 232832 445188
rect 199384 445068 199436 445120
rect 231952 445068 232004 445120
rect 239404 445068 239456 445120
rect 297640 445068 297692 445120
rect 3700 445000 3752 445052
rect 204904 445000 204956 445052
rect 222384 445000 222436 445052
rect 222936 445000 222988 445052
rect 229652 445000 229704 445052
rect 299480 445000 299532 445052
rect 186964 444932 187016 444984
rect 230296 444932 230348 444984
rect 237196 444932 237248 444984
rect 268292 444932 268344 444984
rect 157984 444864 158036 444916
rect 227812 444864 227864 444916
rect 234436 444864 234488 444916
rect 267372 444864 267424 444916
rect 210148 444796 210200 444848
rect 296536 444796 296588 444848
rect 211344 444728 211396 444780
rect 212080 444728 212132 444780
rect 209320 444660 209372 444712
rect 296444 444728 296496 444780
rect 215484 444660 215536 444712
rect 216496 444660 216548 444712
rect 216588 444660 216640 444712
rect 296352 444660 296404 444712
rect 207664 444592 207716 444644
rect 296260 444592 296312 444644
rect 216864 444524 216916 444576
rect 217600 444524 217652 444576
rect 216956 444456 217008 444508
rect 217876 444456 217928 444508
rect 215300 444388 215352 444440
rect 215944 444388 215996 444440
rect 208768 444320 208820 444372
rect 298836 444524 298888 444576
rect 226984 444456 227036 444508
rect 227536 444456 227588 444508
rect 267280 444456 267332 444508
rect 230296 444388 230348 444440
rect 265992 444388 266044 444440
rect 223672 444320 223724 444372
rect 214196 444116 214248 444168
rect 214840 444116 214892 444168
rect 240324 444252 240376 444304
rect 241060 444252 241112 444304
rect 208492 444048 208544 444100
rect 216588 444048 216640 444100
rect 216680 444048 216732 444100
rect 219440 444048 219492 444100
rect 223672 444048 223724 444100
rect 202236 443844 202288 443896
rect 222476 443980 222528 444032
rect 210332 443844 210384 443896
rect 210884 443844 210936 443896
rect 203524 443776 203576 443828
rect 211160 443776 211212 443828
rect 202604 443708 202656 443760
rect 231492 443912 231544 443964
rect 3608 443640 3660 443692
rect 204168 443640 204220 443692
rect 208124 443640 208176 443692
rect 213092 443640 213144 443692
rect 202052 443572 202104 443624
rect 228732 443844 228784 443896
rect 249156 443844 249208 443896
rect 250812 443844 250864 443896
rect 219164 443776 219216 443828
rect 222752 443776 222804 443828
rect 228456 443776 228508 443828
rect 202788 443504 202840 443556
rect 229560 443708 229612 443760
rect 222752 443640 222804 443692
rect 234252 443640 234304 443692
rect 219348 443572 219400 443624
rect 230480 443572 230532 443624
rect 243176 443776 243228 443828
rect 250904 443776 250956 443828
rect 251088 443776 251140 443828
rect 251732 443776 251784 443828
rect 235908 443708 235960 443760
rect 246764 443640 246816 443692
rect 251088 443640 251140 443692
rect 251180 443640 251232 443692
rect 222476 443504 222528 443556
rect 233976 443504 234028 443556
rect 240416 443504 240468 443556
rect 202880 443300 202932 443352
rect 203892 443300 203944 443352
rect 191104 443232 191156 443284
rect 203432 443232 203484 443284
rect 35164 443028 35216 443080
rect 210332 443368 210384 443420
rect 3424 442960 3476 443012
rect 210792 443368 210844 443420
rect 210884 443368 210936 443420
rect 211160 443436 211212 443488
rect 219164 443436 219216 443488
rect 220452 443436 220504 443488
rect 216680 443368 216732 443420
rect 219440 443368 219492 443420
rect 227904 443368 227956 443420
rect 233700 443368 233752 443420
rect 240416 443368 240468 443420
rect 240692 443368 240744 443420
rect 243176 443368 243228 443420
rect 243452 443436 243504 443488
rect 248880 443572 248932 443624
rect 248972 443504 249024 443556
rect 246212 443436 246264 443488
rect 251180 443436 251232 443488
rect 248880 443368 248932 443420
rect 248972 443368 249024 443420
rect 249156 443368 249208 443420
rect 249524 443368 249576 443420
rect 250812 443368 250864 443420
rect 250904 443368 250956 443420
rect 257436 443640 257488 443692
rect 297548 443640 297600 443692
rect 256976 443572 257028 443624
rect 265256 443572 265308 443624
rect 297456 443504 297508 443556
rect 256976 443436 257028 443488
rect 257252 443436 257304 443488
rect 264612 443436 264664 443488
rect 251732 443368 251784 443420
rect 268476 443368 268528 443420
rect 267188 443300 267240 443352
rect 298560 443232 298612 443284
rect 264336 443164 264388 443216
rect 299112 443096 299164 443148
rect 263876 443028 263928 443080
rect 298008 443028 298060 443080
rect 268384 442960 268436 443012
rect 263876 442416 263928 442468
rect 202972 441464 203024 441516
rect 203708 441464 203760 441516
rect 268384 440172 268436 440224
rect 298008 440172 298060 440224
rect 265256 436024 265308 436076
rect 298008 436024 298060 436076
rect 265992 431876 266044 431928
rect 298008 431876 298060 431928
rect 384304 431876 384356 431928
rect 580172 431876 580224 431928
rect 267372 426368 267424 426420
rect 298008 426368 298060 426420
rect 3516 423580 3568 423632
rect 157984 423580 158036 423632
rect 267280 422220 267332 422272
rect 297916 422220 297968 422272
rect 3516 411204 3568 411256
rect 200856 411204 200908 411256
rect 268476 408416 268528 408468
rect 298008 408416 298060 408468
rect 267188 404268 267240 404320
rect 296996 404268 297048 404320
rect 264612 401208 264664 401260
rect 385040 401208 385092 401260
rect 264704 400936 264756 400988
rect 265900 400868 265952 400920
rect 328828 400664 328880 400716
rect 370596 400664 370648 400716
rect 299296 400120 299348 400172
rect 579988 400120 580040 400172
rect 254768 399644 254820 399696
rect 255688 399644 255740 399696
rect 252652 399508 252704 399560
rect 254768 399508 254820 399560
rect 252652 399372 252704 399424
rect 253204 399372 253256 399424
rect 331220 399440 331272 399492
rect 297364 399372 297416 399424
rect 307760 399372 307812 399424
rect 253664 399304 253716 399356
rect 333980 399304 334032 399356
rect 299388 399236 299440 399288
rect 341248 399236 341300 399288
rect 253112 399168 253164 399220
rect 253204 399168 253256 399220
rect 274640 399168 274692 399220
rect 298652 399168 298704 399220
rect 366364 399168 366416 399220
rect 240232 398964 240284 399016
rect 264520 399100 264572 399152
rect 337384 399100 337436 399152
rect 264428 399032 264480 399084
rect 345756 399032 345808 399084
rect 383660 398964 383712 399016
rect 241520 398896 241572 398948
rect 400220 398896 400272 398948
rect 216772 398828 216824 398880
rect 217692 398828 217744 398880
rect 242624 398828 242676 398880
rect 242808 398828 242860 398880
rect 245752 398828 245804 398880
rect 455420 398828 455472 398880
rect 3516 398760 3568 398812
rect 35164 398760 35216 398812
rect 208124 398760 208176 398812
rect 219992 398760 220044 398812
rect 231676 398760 231728 398812
rect 253204 398760 253256 398812
rect 255228 398760 255280 398812
rect 255688 398760 255740 398812
rect 299204 398760 299256 398812
rect 303896 398760 303948 398812
rect 207940 398692 207992 398744
rect 212172 398692 212224 398744
rect 208032 398624 208084 398676
rect 219440 398692 219492 398744
rect 244280 398692 244332 398744
rect 257712 398692 257764 398744
rect 267096 398692 267148 398744
rect 374736 398692 374788 398744
rect 217692 398624 217744 398676
rect 219716 398624 219768 398676
rect 236368 398624 236420 398676
rect 253664 398624 253716 398676
rect 207664 398556 207716 398608
rect 222844 398556 222896 398608
rect 242808 398556 242860 398608
rect 256056 398624 256108 398676
rect 268384 398624 268436 398676
rect 354128 398624 354180 398676
rect 298560 398556 298612 398608
rect 349620 398556 349672 398608
rect 207848 398488 207900 398540
rect 225144 398488 225196 398540
rect 236092 398488 236144 398540
rect 253112 398488 253164 398540
rect 297456 398488 297508 398540
rect 320640 398488 320692 398540
rect 207020 398420 207072 398472
rect 226432 398420 226484 398472
rect 246764 398420 246816 398472
rect 262864 398420 262916 398472
rect 188344 398352 188396 398404
rect 212264 398352 212316 398404
rect 212632 398352 212684 398404
rect 216404 398352 216456 398404
rect 189080 398284 189132 398336
rect 225052 398284 225104 398336
rect 229744 398284 229796 398336
rect 255412 398352 255464 398404
rect 282184 398352 282236 398404
rect 256700 398284 256752 398336
rect 260012 398284 260064 398336
rect 383108 398284 383160 398336
rect 171140 398216 171192 398268
rect 223672 398216 223724 398268
rect 230572 398216 230624 398268
rect 139400 398148 139452 398200
rect 243728 398216 243780 398268
rect 257528 398216 257580 398268
rect 15844 398080 15896 398132
rect 210792 398080 210844 398132
rect 251272 398148 251324 398200
rect 254768 398148 254820 398200
rect 543740 398148 543792 398200
rect 221188 398080 221240 398132
rect 242072 398080 242124 398132
rect 209780 398012 209832 398064
rect 212632 398012 212684 398064
rect 216312 398012 216364 398064
rect 223120 398012 223172 398064
rect 254032 398080 254084 398132
rect 561680 398080 561732 398132
rect 256148 398012 256200 398064
rect 212172 397944 212224 397996
rect 218888 397944 218940 397996
rect 209136 397876 209188 397928
rect 217784 397876 217836 397928
rect 246212 397876 246264 397928
rect 260196 397944 260248 397996
rect 254032 397876 254084 397928
rect 260104 397876 260156 397928
rect 215300 397808 215352 397860
rect 223028 397808 223080 397860
rect 232596 397808 232648 397860
rect 209228 397672 209280 397724
rect 218336 397672 218388 397724
rect 219992 397672 220044 397724
rect 227444 397672 227496 397724
rect 210332 397604 210384 397656
rect 215852 397604 215904 397656
rect 219624 397604 219676 397656
rect 220360 397604 220412 397656
rect 220820 397604 220872 397656
rect 227352 397604 227404 397656
rect 238760 397808 238812 397860
rect 242808 397808 242860 397860
rect 245660 397808 245712 397860
rect 239312 397740 239364 397792
rect 246764 397740 246816 397792
rect 240416 397672 240468 397724
rect 246212 397672 246264 397724
rect 253112 397808 253164 397860
rect 251272 397740 251324 397792
rect 259460 397740 259512 397792
rect 254032 397672 254084 397724
rect 239680 397604 239732 397656
rect 239864 397604 239916 397656
rect 243912 397604 243964 397656
rect 244832 397604 244884 397656
rect 258724 397672 258776 397724
rect 212908 397536 212960 397588
rect 213460 397536 213512 397588
rect 213920 397536 213972 397588
rect 217232 397536 217284 397588
rect 209320 397468 209372 397520
rect 210792 397468 210844 397520
rect 212172 397468 212224 397520
rect 213828 397468 213880 397520
rect 222200 397536 222252 397588
rect 227168 397536 227220 397588
rect 234712 397536 234764 397588
rect 240048 397536 240100 397588
rect 240968 397536 241020 397588
rect 246948 397536 247000 397588
rect 212908 397400 212960 397452
rect 220360 397468 220412 397520
rect 220912 397468 220964 397520
rect 222384 397468 222436 397520
rect 226432 397468 226484 397520
rect 227812 397468 227864 397520
rect 238208 397468 238260 397520
rect 242532 397468 242584 397520
rect 243176 397468 243228 397520
rect 257436 397604 257488 397656
rect 525800 397604 525852 397656
rect 254308 397536 254360 397588
rect 564440 397536 564492 397588
rect 256792 397468 256844 397520
rect 582380 397468 582432 397520
rect 237472 397400 237524 397452
rect 238392 397400 238444 397452
rect 210792 397332 210844 397384
rect 224684 397332 224736 397384
rect 37280 397264 37332 397316
rect 213276 397264 213328 397316
rect 245936 397264 245988 397316
rect 257344 397264 257396 397316
rect 212540 397196 212592 397248
rect 213368 397196 213420 397248
rect 198740 397128 198792 397180
rect 225788 397128 225840 397180
rect 234252 397128 234304 397180
rect 162860 397060 162912 397112
rect 215300 397060 215352 397112
rect 151820 396992 151872 397044
rect 212908 396992 212960 397044
rect 213000 396992 213052 397044
rect 213368 396992 213420 397044
rect 214104 396992 214156 397044
rect 214564 396992 214616 397044
rect 218060 396992 218112 397044
rect 218888 396992 218940 397044
rect 144920 396924 144972 396976
rect 221648 396924 221700 396976
rect 131120 396856 131172 396908
rect 40040 396788 40092 396840
rect 212540 396788 212592 396840
rect 210148 396720 210200 396772
rect 210608 396720 210660 396772
rect 211252 396720 211304 396772
rect 211988 396720 212040 396772
rect 212724 396720 212776 396772
rect 213736 396720 213788 396772
rect 209872 396652 209924 396704
rect 210424 396652 210476 396704
rect 211620 396652 211672 396704
rect 211896 396652 211948 396704
rect 213000 396652 213052 396704
rect 213644 396652 213696 396704
rect 218152 396856 218204 396908
rect 218796 396856 218848 396908
rect 219440 396856 219492 396908
rect 220084 396856 220136 396908
rect 222384 396856 222436 396908
rect 222660 396856 222712 396908
rect 237380 397128 237432 397180
rect 237932 397128 237984 397180
rect 237656 396992 237708 397044
rect 237932 396992 237984 397044
rect 307760 396856 307812 396908
rect 215300 396788 215352 396840
rect 215484 396720 215536 396772
rect 215944 396720 215996 396772
rect 218428 396720 218480 396772
rect 218612 396720 218664 396772
rect 219716 396788 219768 396840
rect 220176 396788 220228 396840
rect 222568 396788 222620 396840
rect 222844 396788 222896 396840
rect 223856 396788 223908 396840
rect 224316 396788 224368 396840
rect 236736 396788 236788 396840
rect 339500 396788 339552 396840
rect 223396 396720 223448 396772
rect 241152 396720 241204 396772
rect 396080 396720 396132 396772
rect 220544 396652 220596 396704
rect 221096 396652 221148 396704
rect 221556 396652 221608 396704
rect 224316 396652 224368 396704
rect 224776 396652 224828 396704
rect 210516 396584 210568 396636
rect 211344 396584 211396 396636
rect 212080 396584 212132 396636
rect 212908 396584 212960 396636
rect 213552 396584 213604 396636
rect 214196 396584 214248 396636
rect 215116 396584 215168 396636
rect 215760 396584 215812 396636
rect 216496 396584 216548 396636
rect 218244 396584 218296 396636
rect 219256 396584 219308 396636
rect 219808 396584 219860 396636
rect 220452 396584 220504 396636
rect 221004 396584 221056 396636
rect 221832 396584 221884 396636
rect 223764 396584 223816 396636
rect 224868 396584 224920 396636
rect 232504 396584 232556 396636
rect 209964 396516 210016 396568
rect 210056 396516 210108 396568
rect 210976 396516 211028 396568
rect 211436 396516 211488 396568
rect 212448 396516 212500 396568
rect 214380 396516 214432 396568
rect 215208 396516 215260 396568
rect 215576 396516 215628 396568
rect 216588 396516 216640 396568
rect 216864 396516 216916 396568
rect 217876 396516 217928 396568
rect 218336 396516 218388 396568
rect 218796 396516 218848 396568
rect 219624 396516 219676 396568
rect 220636 396516 220688 396568
rect 221280 396516 221332 396568
rect 221924 396516 221976 396568
rect 222476 396516 222528 396568
rect 223304 396516 223356 396568
rect 224040 396516 224092 396568
rect 224408 396516 224460 396568
rect 242164 396584 242216 396636
rect 213920 396448 213972 396500
rect 215024 396448 215076 396500
rect 218704 396448 218756 396500
rect 219164 396448 219216 396500
rect 219900 396448 219952 396500
rect 220268 396448 220320 396500
rect 221372 396448 221424 396500
rect 222108 396448 222160 396500
rect 232688 396448 232740 396500
rect 209780 396380 209832 396432
rect 210608 396380 210660 396432
rect 213184 396380 213236 396432
rect 215300 396380 215352 396432
rect 217048 396380 217100 396432
rect 217600 396380 217652 396432
rect 218520 396380 218572 396432
rect 219072 396380 219124 396432
rect 242348 396380 242400 396432
rect 215668 396312 215720 396364
rect 216128 396312 216180 396364
rect 217232 396312 217284 396364
rect 217968 396312 218020 396364
rect 218336 396312 218388 396364
rect 218980 396312 219032 396364
rect 217140 396244 217192 396296
rect 217416 396244 217468 396296
rect 219992 396176 220044 396228
rect 220728 396176 220780 396228
rect 220912 396176 220964 396228
rect 222016 396176 222068 396228
rect 244188 396108 244240 396160
rect 245384 396108 245436 396160
rect 210424 396040 210476 396092
rect 210792 396040 210844 396092
rect 210240 395972 210292 396024
rect 211068 395972 211120 396024
rect 217324 395972 217376 396024
rect 217692 395972 217744 396024
rect 220084 395972 220136 396024
rect 226892 395972 226944 396024
rect 204904 395836 204956 395888
rect 224132 395836 224184 395888
rect 230848 395836 230900 395888
rect 231492 395836 231544 395888
rect 115940 395564 115992 395616
rect 218060 395768 218112 395820
rect 231952 395768 232004 395820
rect 232872 395768 232924 395820
rect 109040 395496 109092 395548
rect 218152 395700 218204 395752
rect 246764 395700 246816 395752
rect 372620 395700 372672 395752
rect 215944 395632 215996 395684
rect 216312 395632 216364 395684
rect 247684 395632 247736 395684
rect 248052 395632 248104 395684
rect 249248 395632 249300 395684
rect 499580 395632 499632 395684
rect 214472 395564 214524 395616
rect 214656 395564 214708 395616
rect 250352 395564 250404 395616
rect 514760 395564 514812 395616
rect 93860 395428 93912 395480
rect 216680 395496 216732 395548
rect 251456 395496 251508 395548
rect 528560 395496 528612 395548
rect 214472 395428 214524 395480
rect 214932 395428 214984 395480
rect 252008 395428 252060 395480
rect 535460 395428 535512 395480
rect 86960 395360 87012 395412
rect 214748 395360 214800 395412
rect 253204 395360 253256 395412
rect 549260 395360 549312 395412
rect 77300 395292 77352 395344
rect 216404 395292 216456 395344
rect 255228 395292 255280 395344
rect 571340 395292 571392 395344
rect 240324 395088 240376 395140
rect 240968 395088 241020 395140
rect 242992 395088 243044 395140
rect 243728 395088 243780 395140
rect 248696 395020 248748 395072
rect 249248 395020 249300 395072
rect 214012 394952 214064 395004
rect 214840 394952 214892 395004
rect 213276 394884 213328 394936
rect 213828 394884 213880 394936
rect 253940 394748 253992 394800
rect 254768 394748 254820 394800
rect 236000 394612 236052 394664
rect 244188 394612 244240 394664
rect 244556 394612 244608 394664
rect 244832 394612 244884 394664
rect 247040 394612 247092 394664
rect 236828 394544 236880 394596
rect 244096 394544 244148 394596
rect 244372 394544 244424 394596
rect 244924 394544 244976 394596
rect 249892 394544 249944 394596
rect 250260 394544 250312 394596
rect 251548 394612 251600 394664
rect 252192 394612 252244 394664
rect 253940 394612 253992 394664
rect 254584 394612 254636 394664
rect 255964 394544 256016 394596
rect 237472 394476 237524 394528
rect 244004 394476 244056 394528
rect 244280 394476 244332 394528
rect 244648 394476 244700 394528
rect 245752 394476 245804 394528
rect 246028 394476 246080 394528
rect 250168 394476 250220 394528
rect 250812 394476 250864 394528
rect 251548 394476 251600 394528
rect 251916 394476 251968 394528
rect 252836 394476 252888 394528
rect 253204 394476 253256 394528
rect 254124 394476 254176 394528
rect 254400 394476 254452 394528
rect 227260 394408 227312 394460
rect 234344 394408 234396 394460
rect 307852 394408 307904 394460
rect 209044 394204 209096 394256
rect 219440 394204 219492 394256
rect 195980 394136 196032 394188
rect 225604 394204 225656 394256
rect 235172 394340 235224 394392
rect 228456 394272 228508 394324
rect 228732 394272 228784 394324
rect 233792 394272 233844 394324
rect 234068 394272 234120 394324
rect 234712 394272 234764 394324
rect 235264 394272 235316 394324
rect 227352 394204 227404 394256
rect 240140 394272 240192 394324
rect 241152 394272 241204 394324
rect 241520 394272 241572 394324
rect 241796 394272 241848 394324
rect 242900 394272 242952 394324
rect 243176 394272 243228 394324
rect 224132 394136 224184 394188
rect 224500 394136 224552 394188
rect 231952 394136 232004 394188
rect 232228 394136 232280 394188
rect 234620 394136 234672 394188
rect 235172 394136 235224 394188
rect 239036 394136 239088 394188
rect 168380 394068 168432 394120
rect 223488 394068 223540 394120
rect 232412 394068 232464 394120
rect 232596 394068 232648 394120
rect 234988 394068 235040 394120
rect 235356 394068 235408 394120
rect 241704 394136 241756 394188
rect 242164 394136 242216 394188
rect 242808 394204 242860 394256
rect 243544 394204 243596 394256
rect 318800 394340 318852 394392
rect 244188 394272 244240 394324
rect 329840 394272 329892 394324
rect 244096 394204 244148 394256
rect 340880 394204 340932 394256
rect 244004 394136 244056 394188
rect 347780 394136 347832 394188
rect 143540 394000 143592 394052
rect 221464 394000 221516 394052
rect 228548 394000 228600 394052
rect 234620 394000 234672 394052
rect 236000 394000 236052 394052
rect 236920 394000 236972 394052
rect 241980 394000 242032 394052
rect 242256 394000 242308 394052
rect 242716 394068 242768 394120
rect 365720 394068 365772 394120
rect 368480 394000 368532 394052
rect 63500 393932 63552 393984
rect 212448 393932 212500 393984
rect 219440 393932 219492 393984
rect 220176 393932 220228 393984
rect 225604 393932 225656 393984
rect 226248 393932 226300 393984
rect 226616 393932 226668 393984
rect 226984 393932 227036 393984
rect 227812 393932 227864 393984
rect 227996 393932 228048 393984
rect 228088 393932 228140 393984
rect 228824 393932 228876 393984
rect 229284 393932 229336 393984
rect 230112 393932 230164 393984
rect 230756 393932 230808 393984
rect 230940 393932 230992 393984
rect 231860 393932 231912 393984
rect 232412 393932 232464 393984
rect 233516 393932 233568 393984
rect 233792 393932 233844 393984
rect 236092 393932 236144 393984
rect 236644 393932 236696 393984
rect 237472 393932 237524 393984
rect 238024 393932 238076 393984
rect 238760 393932 238812 393984
rect 239404 393932 239456 393984
rect 240416 393932 240468 393984
rect 240876 393932 240928 393984
rect 241796 393932 241848 393984
rect 242348 393932 242400 393984
rect 242992 393932 243044 393984
rect 243268 393932 243320 393984
rect 243912 393932 243964 393984
rect 379520 393932 379572 393984
rect 225144 393864 225196 393916
rect 225696 393864 225748 393916
rect 229376 393864 229428 393916
rect 234160 393864 234212 393916
rect 235264 393864 235316 393916
rect 240232 393864 240284 393916
rect 240784 393864 240836 393916
rect 245660 393864 245712 393916
rect 246304 393864 246356 393916
rect 247224 393864 247276 393916
rect 225512 393796 225564 393848
rect 226156 393796 226208 393848
rect 229284 393796 229336 393848
rect 229560 393796 229612 393848
rect 230572 393796 230624 393848
rect 231124 393796 231176 393848
rect 231860 393796 231912 393848
rect 232688 393796 232740 393848
rect 233240 393796 233292 393848
rect 233516 393796 233568 393848
rect 225236 393728 225288 393780
rect 226064 393728 226116 393780
rect 230664 393728 230716 393780
rect 231400 393728 231452 393780
rect 232044 393728 232096 393780
rect 232780 393728 232832 393780
rect 238852 393796 238904 393848
rect 239128 393796 239180 393848
rect 240324 393796 240376 393848
rect 241060 393796 241112 393848
rect 241612 393796 241664 393848
rect 242440 393796 242492 393848
rect 243084 393796 243136 393848
rect 243452 393796 243504 393848
rect 245844 393796 245896 393848
rect 246580 393796 246632 393848
rect 243268 393728 243320 393780
rect 243636 393728 243688 393780
rect 245936 393728 245988 393780
rect 246120 393728 246172 393780
rect 248420 393864 248472 393916
rect 248788 393864 248840 393916
rect 249800 393864 249852 393916
rect 250168 393864 250220 393916
rect 250260 393864 250312 393916
rect 250628 393864 250680 393916
rect 251732 393864 251784 393916
rect 251916 393864 251968 393916
rect 254584 393864 254636 393916
rect 254952 393864 255004 393916
rect 251364 393796 251416 393848
rect 251640 393796 251692 393848
rect 252652 393796 252704 393848
rect 252836 393796 252888 393848
rect 253020 393796 253072 393848
rect 253388 393796 253440 393848
rect 254308 393796 254360 393848
rect 254492 393796 254544 393848
rect 255320 393796 255372 393848
rect 255596 393796 255648 393848
rect 248420 393728 248472 393780
rect 249340 393728 249392 393780
rect 251272 393728 251324 393780
rect 252100 393728 252152 393780
rect 254216 393728 254268 393780
rect 254676 393728 254728 393780
rect 226432 393660 226484 393712
rect 227076 393660 227128 393712
rect 227996 393660 228048 393712
rect 228364 393660 228416 393712
rect 230848 393660 230900 393712
rect 231216 393660 231268 393712
rect 234896 393660 234948 393712
rect 235080 393660 235132 393712
rect 235448 393660 235500 393712
rect 243084 393660 243136 393712
rect 243820 393660 243872 393712
rect 244372 393660 244424 393712
rect 245200 393660 245252 393712
rect 247408 393660 247460 393712
rect 248696 393660 248748 393712
rect 249156 393660 249208 393712
rect 252468 393660 252520 393712
rect 253112 393660 253164 393712
rect 254032 393660 254084 393712
rect 254492 393660 254544 393712
rect 226892 393592 226944 393644
rect 227628 393592 227680 393644
rect 227720 393592 227772 393644
rect 228088 393592 228140 393644
rect 246120 393592 246172 393644
rect 246396 393592 246448 393644
rect 227904 393524 227956 393576
rect 228456 393524 228508 393576
rect 230388 393524 230440 393576
rect 231216 393524 231268 393576
rect 239128 393524 239180 393576
rect 239588 393524 239640 393576
rect 254032 393524 254084 393576
rect 254860 393524 254912 393576
rect 236276 393456 236328 393508
rect 236460 393456 236512 393508
rect 239036 393456 239088 393508
rect 239496 393456 239548 393508
rect 231492 392844 231544 392896
rect 257620 392844 257672 392896
rect 232872 392776 232924 392828
rect 277400 392776 277452 392828
rect 238392 392708 238444 392760
rect 349160 392708 349212 392760
rect 164240 392640 164292 392692
rect 215944 392640 215996 392692
rect 245016 392640 245068 392692
rect 445760 392640 445812 392692
rect 34520 392572 34572 392624
rect 213368 392572 213420 392624
rect 248052 392572 248104 392624
rect 480260 392572 480312 392624
rect 249984 392300 250036 392352
rect 250536 392300 250588 392352
rect 251180 392300 251232 392352
rect 251824 392300 251876 392352
rect 229192 392164 229244 392216
rect 229468 392164 229520 392216
rect 233424 392164 233476 392216
rect 233700 392164 233752 392216
rect 237564 392164 237616 392216
rect 237748 392164 237800 392216
rect 233332 392096 233384 392148
rect 233884 392096 233936 392148
rect 229100 392028 229152 392080
rect 229744 392028 229796 392080
rect 237564 392028 237616 392080
rect 238300 392028 238352 392080
rect 229284 391892 229336 391944
rect 230020 391892 230072 391944
rect 228732 391824 228784 391876
rect 233516 391824 233568 391876
rect 225420 391688 225472 391740
rect 225972 391688 226024 391740
rect 240048 391484 240100 391536
rect 313280 391484 313332 391536
rect 240968 391416 241020 391468
rect 385040 391416 385092 391468
rect 243728 391348 243780 391400
rect 419540 391348 419592 391400
rect 236368 391280 236420 391332
rect 184940 391212 184992 391264
rect 224316 391212 224368 391264
rect 245384 391280 245436 391332
rect 437480 391280 437532 391332
rect 249248 391212 249300 391264
rect 492680 391212 492732 391264
rect 236460 391076 236512 391128
rect 252836 391008 252888 391060
rect 253296 391008 253348 391060
rect 247316 390396 247368 390448
rect 247776 390396 247828 390448
rect 247592 390328 247644 390380
rect 247776 390124 247828 390176
rect 234068 389784 234120 389836
rect 300860 389784 300912 389836
rect 233516 389376 233568 389428
rect 233976 389376 234028 389428
rect 233424 389240 233476 389292
rect 233792 389172 233844 389224
rect 233884 389172 233936 389224
rect 234160 389172 234212 389224
rect 227168 386520 227220 386572
rect 227536 386520 227588 386572
rect 299112 379448 299164 379500
rect 580172 379448 580224 379500
rect 3056 372512 3108 372564
rect 106924 372512 106976 372564
rect 296628 365644 296680 365696
rect 580172 365644 580224 365696
rect 3516 358708 3568 358760
rect 184204 358708 184256 358760
rect 23480 358028 23532 358080
rect 208216 358028 208268 358080
rect 237932 356668 237984 356720
rect 350540 356668 350592 356720
rect 235264 355648 235316 355700
rect 316040 355648 316092 355700
rect 235448 355580 235500 355632
rect 324412 355580 324464 355632
rect 113180 355512 113232 355564
rect 218704 355512 218756 355564
rect 242440 355512 242492 355564
rect 357440 355512 357492 355564
rect 88340 355444 88392 355496
rect 213276 355444 213328 355496
rect 239220 355444 239272 355496
rect 367100 355444 367152 355496
rect 73160 355376 73212 355428
rect 215852 355376 215904 355428
rect 239312 355376 239364 355428
rect 371240 355376 371292 355428
rect 45560 355308 45612 355360
rect 204996 355308 205048 355360
rect 246672 355308 246724 355360
rect 393320 355308 393372 355360
rect 78680 354356 78732 354408
rect 215760 354356 215812 354408
rect 56600 354288 56652 354340
rect 211896 354288 211948 354340
rect 231308 354288 231360 354340
rect 269120 354288 269172 354340
rect 42800 354220 42852 354272
rect 213000 354220 213052 354272
rect 232596 354220 232648 354272
rect 284300 354220 284352 354272
rect 41420 354152 41472 354204
rect 212908 354152 212960 354204
rect 238024 354152 238076 354204
rect 357532 354152 357584 354204
rect 19340 354084 19392 354136
rect 211620 354084 211672 354136
rect 240784 354084 240836 354136
rect 397460 354084 397512 354136
rect 19432 354016 19484 354068
rect 211712 354016 211764 354068
rect 229744 354016 229796 354068
rect 242072 354016 242124 354068
rect 251916 354016 251968 354068
rect 531320 354016 531372 354068
rect 13820 353948 13872 354000
rect 210700 353948 210752 354000
rect 229836 353948 229888 354000
rect 251640 353948 251692 354000
rect 254676 353948 254728 354000
rect 560300 353948 560352 354000
rect 231216 352792 231268 352844
rect 259552 352792 259604 352844
rect 157340 352724 157392 352776
rect 222752 352724 222804 352776
rect 231032 352724 231084 352776
rect 266360 352724 266412 352776
rect 104900 352656 104952 352708
rect 218612 352656 218664 352708
rect 257712 352656 257764 352708
rect 436100 352656 436152 352708
rect 52460 352588 52512 352640
rect 214656 352588 214708 352640
rect 250536 352588 250588 352640
rect 512000 352588 512052 352640
rect 3516 352520 3568 352572
rect 201960 352520 202012 352572
rect 213276 352520 213328 352572
rect 227076 352520 227128 352572
rect 228364 352520 228416 352572
rect 235264 352520 235316 352572
rect 251824 352520 251876 352572
rect 524420 352520 524472 352572
rect 204260 351364 204312 351416
rect 225604 351364 225656 351416
rect 182180 351296 182232 351348
rect 224132 351296 224184 351348
rect 151912 351228 151964 351280
rect 221372 351228 221424 351280
rect 236552 351228 236604 351280
rect 342260 351228 342312 351280
rect 4160 351160 4212 351212
rect 209320 351160 209372 351212
rect 253296 351160 253348 351212
rect 554780 351160 554832 351212
rect 222752 350548 222804 350600
rect 226892 350548 226944 350600
rect 254584 347012 254636 347064
rect 572720 347012 572772 347064
rect 3148 346332 3200 346384
rect 202052 346332 202104 346384
rect 260196 335996 260248 336048
rect 460940 335996 460992 336048
rect 299020 325592 299072 325644
rect 579896 325592 579948 325644
rect 2780 320084 2832 320136
rect 6276 320084 6328 320136
rect 296536 313216 296588 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 14464 306280 14516 306332
rect 258816 302880 258868 302932
rect 449900 302880 449952 302932
rect 3240 293904 3292 293956
rect 202788 293904 202840 293956
rect 298928 273164 298980 273216
rect 579896 273164 579948 273216
rect 3240 267656 3292 267708
rect 186964 267656 187016 267708
rect 296444 259360 296496 259412
rect 579804 259360 579856 259412
rect 3148 254736 3200 254788
rect 6184 254736 6236 254788
rect 298836 245556 298888 245608
rect 580172 245556 580224 245608
rect 3332 241408 3384 241460
rect 191104 241408 191156 241460
rect 265808 233180 265860 233232
rect 580172 233180 580224 233232
rect 246304 228352 246356 228404
rect 386420 228352 386472 228404
rect 296352 219376 296404 219428
rect 579896 219376 579948 219428
rect 3148 215228 3200 215280
rect 203616 215228 203668 215280
rect 264336 206932 264388 206984
rect 580172 206932 580224 206984
rect 3332 202784 3384 202836
rect 202604 202784 202656 202836
rect 298744 193128 298796 193180
rect 580172 193128 580224 193180
rect 262864 182792 262916 182844
rect 467840 182792 467892 182844
rect 296260 179324 296312 179376
rect 579988 179324 580040 179376
rect 233792 177692 233844 177744
rect 293960 177692 294012 177744
rect 233976 177624 234028 177676
rect 298100 177624 298152 177676
rect 203064 177556 203116 177608
rect 225512 177556 225564 177608
rect 240692 177556 240744 177608
rect 382280 177556 382332 177608
rect 201500 177488 201552 177540
rect 225420 177488 225472 177540
rect 240600 177488 240652 177540
rect 390560 177488 390612 177540
rect 133880 177420 133932 177472
rect 219992 177420 220044 177472
rect 247684 177420 247736 177472
rect 478880 177420 478932 177472
rect 126980 177352 127032 177404
rect 219900 177352 219952 177404
rect 250444 177352 250496 177404
rect 518900 177352 518952 177404
rect 77392 177284 77444 177336
rect 210608 177284 210660 177336
rect 215760 177284 215812 177336
rect 226800 177284 226852 177336
rect 251732 177284 251784 177336
rect 532700 177284 532752 177336
rect 38660 175924 38712 175976
rect 206468 175924 206520 175976
rect 102140 171776 102192 171828
rect 209228 171776 209280 171828
rect 272524 166948 272576 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 199384 164160 199436 164212
rect 3332 150356 3384 150408
rect 202696 150356 202748 150408
rect 296076 139340 296128 139392
rect 580172 139340 580224 139392
rect 267004 126896 267056 126948
rect 580172 126896 580224 126948
rect 265716 113092 265768 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 200764 111732 200816 111784
rect 296168 100648 296220 100700
rect 580172 100648 580224 100700
rect 3240 97928 3292 97980
rect 202512 97928 202564 97980
rect 249064 88952 249116 89004
rect 502340 88952 502392 89004
rect 235356 87728 235408 87780
rect 316132 87728 316184 87780
rect 242256 87660 242308 87712
rect 407120 87660 407172 87712
rect 244924 87592 244976 87644
rect 448520 87592 448572 87644
rect 264244 86912 264296 86964
rect 580172 86912 580224 86964
rect 247592 86300 247644 86352
rect 481640 86300 481692 86352
rect 250352 86232 250404 86284
rect 514852 86232 514904 86284
rect 3332 85484 3384 85536
rect 202420 85484 202472 85536
rect 239404 84872 239456 84924
rect 285680 84872 285732 84924
rect 254492 84804 254544 84856
rect 563060 84804 563112 84856
rect 242164 83444 242216 83496
rect 402980 83444 403032 83496
rect 230940 82152 230992 82204
rect 262220 82152 262272 82204
rect 247500 82084 247552 82136
rect 477500 82084 477552 82136
rect 265624 73108 265676 73160
rect 580172 73108 580224 73160
rect 3332 71680 3384 71732
rect 202328 71680 202380 71732
rect 295984 60664 296036 60716
rect 580172 60664 580224 60716
rect 3332 59304 3384 59356
rect 202236 59304 202288 59356
rect 202972 58624 203024 58676
rect 580264 58624 580316 58676
rect 260104 48968 260156 49020
rect 454040 48968 454092 49020
rect 211620 46248 211672 46300
rect 226708 46248 226760 46300
rect 160100 46180 160152 46232
rect 222660 46180 222712 46232
rect 124220 37884 124272 37936
rect 208124 37884 208176 37936
rect 95240 35164 95292 35216
rect 209136 35164 209188 35216
rect 258724 35164 258776 35216
rect 443000 35164 443052 35216
rect 202880 33056 202932 33108
rect 580172 33056 580224 33108
rect 3424 32988 3476 33040
rect 203524 32988 203576 33040
rect 256240 28296 256292 28348
rect 494060 28296 494112 28348
rect 248972 28228 249024 28280
rect 498200 28228 498252 28280
rect 256148 26936 256200 26988
rect 407212 26936 407264 26988
rect 256056 26868 256108 26920
rect 415400 26868 415452 26920
rect 232504 25984 232556 26036
rect 287060 25984 287112 26036
rect 235172 25916 235224 25968
rect 311900 25916 311952 25968
rect 235080 25848 235132 25900
rect 322940 25848 322992 25900
rect 236460 25780 236512 25832
rect 332600 25780 332652 25832
rect 239128 25712 239180 25764
rect 375380 25712 375432 25764
rect 243544 25644 243596 25696
rect 425060 25644 425112 25696
rect 244740 25576 244792 25628
rect 440240 25576 440292 25628
rect 244832 25508 244884 25560
rect 447140 25508 447192 25560
rect 232412 24488 232464 24540
rect 276020 24488 276072 24540
rect 232320 24420 232372 24472
rect 280160 24420 280212 24472
rect 250260 24352 250312 24404
rect 517520 24352 517572 24404
rect 253112 24284 253164 24336
rect 542360 24284 542412 24336
rect 253204 24216 253256 24268
rect 546500 24216 546552 24268
rect 253020 24148 253072 24200
rect 553400 24148 553452 24200
rect 254400 24080 254452 24132
rect 564532 24080 564584 24132
rect 236368 23128 236420 23180
rect 336740 23128 336792 23180
rect 246120 23060 246172 23112
rect 463700 23060 463752 23112
rect 247408 22992 247460 23044
rect 473360 22992 473412 23044
rect 248788 22924 248840 22976
rect 490012 22924 490064 22976
rect 248880 22856 248932 22908
rect 496820 22856 496872 22908
rect 250168 22788 250220 22840
rect 506572 22788 506624 22840
rect 5540 22720 5592 22772
rect 15844 22720 15896 22772
rect 250076 22720 250128 22772
rect 510620 22720 510672 22772
rect 241980 21836 242032 21888
rect 409880 21836 409932 21888
rect 243452 21768 243504 21820
rect 420920 21768 420972 21820
rect 243360 21700 243412 21752
rect 423680 21700 423732 21752
rect 243268 21632 243320 21684
rect 427820 21632 427872 21684
rect 244556 21564 244608 21616
rect 438860 21564 438912 21616
rect 244648 21496 244700 21548
rect 441620 21496 441672 21548
rect 246028 21428 246080 21480
rect 456892 21428 456944 21480
rect 245936 21360 245988 21412
rect 459560 21360 459612 21412
rect 3424 20612 3476 20664
rect 202144 20612 202196 20664
rect 237748 20204 237800 20256
rect 349252 20204 349304 20256
rect 237840 20136 237892 20188
rect 353300 20136 353352 20188
rect 239036 20068 239088 20120
rect 374000 20068 374052 20120
rect 240508 20000 240560 20052
rect 389180 20000 389232 20052
rect 240416 19932 240468 19984
rect 391940 19932 391992 19984
rect 233700 19048 233752 19100
rect 296720 19048 296772 19100
rect 233608 18980 233660 19032
rect 299480 18980 299532 19032
rect 233516 18912 233568 18964
rect 303620 18912 303672 18964
rect 234804 18844 234856 18896
rect 314660 18844 314712 18896
rect 234988 18776 235040 18828
rect 317420 18776 317472 18828
rect 234896 18708 234948 18760
rect 321560 18708 321612 18760
rect 236184 18640 236236 18692
rect 332692 18640 332744 18692
rect 236276 18572 236328 18624
rect 335360 18572 335412 18624
rect 232136 17620 232188 17672
rect 278780 17620 278832 17672
rect 232228 17552 232280 17604
rect 282920 17552 282972 17604
rect 251548 17484 251600 17536
rect 534080 17484 534132 17536
rect 252744 17416 252796 17468
rect 545120 17416 545172 17468
rect 252928 17348 252980 17400
rect 547880 17348 547932 17400
rect 252836 17280 252888 17332
rect 552020 17280 552072 17332
rect 180800 17212 180852 17264
rect 224040 17212 224092 17264
rect 254308 17212 254360 17264
rect 567200 17212 567252 17264
rect 243176 16260 243228 16312
rect 418528 16260 418580 16312
rect 248696 16192 248748 16244
rect 498936 16192 498988 16244
rect 249892 16124 249944 16176
rect 509608 16124 509660 16176
rect 136456 16056 136508 16108
rect 220176 16056 220228 16108
rect 249800 16056 249852 16108
rect 513380 16056 513432 16108
rect 71504 15988 71556 16040
rect 210516 15988 210568 16040
rect 249984 15988 250036 16040
rect 517152 15988 517204 16040
rect 35992 15920 36044 15972
rect 212816 15920 212868 15972
rect 251456 15920 251508 15972
rect 527824 15920 527876 15972
rect 9680 15852 9732 15904
rect 210240 15852 210292 15904
rect 251364 15852 251416 15904
rect 531412 15852 531464 15904
rect 163504 14968 163556 15020
rect 218428 14968 218480 15020
rect 112352 14900 112404 14952
rect 218520 14900 218572 14952
rect 98184 14832 98236 14884
rect 217232 14832 217284 14884
rect 91560 14764 91612 14816
rect 217140 14764 217192 14816
rect 247132 14764 247184 14816
rect 473452 14764 473504 14816
rect 75000 14696 75052 14748
rect 215668 14696 215720 14748
rect 247224 14696 247276 14748
rect 476488 14696 476540 14748
rect 44180 14628 44232 14680
rect 211804 14628 211856 14680
rect 247316 14628 247368 14680
rect 481732 14628 481784 14680
rect 27712 14560 27764 14612
rect 211436 14560 211488 14612
rect 248512 14560 248564 14612
rect 492312 14560 492364 14612
rect 22560 14492 22612 14544
rect 211344 14492 211396 14544
rect 248604 14492 248656 14544
rect 495440 14492 495492 14544
rect 17960 14424 18012 14476
rect 211528 14424 211580 14476
rect 254216 14424 254268 14476
rect 570328 14424 570380 14476
rect 80888 13472 80940 13524
rect 215576 13472 215628 13524
rect 243084 13472 243136 13524
rect 430856 13472 430908 13524
rect 63224 13404 63276 13456
rect 214380 13404 214432 13456
rect 244280 13404 244332 13456
rect 440332 13404 440384 13456
rect 59360 13336 59412 13388
rect 214472 13336 214524 13388
rect 244464 13336 244516 13388
rect 445024 13336 445076 13388
rect 56048 13268 56100 13320
rect 214564 13268 214616 13320
rect 244372 13268 244424 13320
rect 448612 13268 448664 13320
rect 52552 13200 52604 13252
rect 214288 13200 214340 13252
rect 245752 13200 245804 13252
rect 459192 13200 459244 13252
rect 8760 13132 8812 13184
rect 210056 13132 210108 13184
rect 245660 13132 245712 13184
rect 462320 13132 462372 13184
rect 3424 13064 3476 13116
rect 210148 13064 210200 13116
rect 245844 13064 245896 13116
rect 465816 13064 465868 13116
rect 114744 12180 114796 12232
rect 218244 12180 218296 12232
rect 110420 12112 110472 12164
rect 218336 12112 218388 12164
rect 108120 12044 108172 12096
rect 218888 12044 218940 12096
rect 240324 12044 240376 12096
rect 395344 12044 395396 12096
rect 44272 11976 44324 12028
rect 212724 11976 212776 12028
rect 241704 11976 241756 12028
rect 402520 11976 402572 12028
rect 36728 11908 36780 11960
rect 213092 11908 213144 11960
rect 241888 11908 241940 11960
rect 406016 11908 406068 11960
rect 33600 11840 33652 11892
rect 213460 11840 213512 11892
rect 241796 11840 241848 11892
rect 409144 11840 409196 11892
rect 26240 11772 26292 11824
rect 212356 11772 212408 11824
rect 242992 11772 243044 11824
rect 423772 11772 423824 11824
rect 21824 11704 21876 11756
rect 211252 11704 211304 11756
rect 242900 11704 242952 11756
rect 426808 11704 426860 11756
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 159364 10752 159416 10804
rect 218796 10752 218848 10804
rect 97448 10684 97500 10736
rect 216864 10684 216916 10736
rect 93952 10616 94004 10668
rect 217048 10616 217100 10668
rect 238944 10616 238996 10668
rect 365812 10616 365864 10668
rect 89904 10548 89956 10600
rect 216956 10548 217008 10600
rect 238852 10548 238904 10600
rect 370136 10548 370188 10600
rect 86408 10480 86460 10532
rect 216772 10480 216824 10532
rect 238760 10480 238812 10532
rect 374092 10480 374144 10532
rect 75920 10412 75972 10464
rect 216128 10412 216180 10464
rect 240140 10412 240192 10464
rect 387800 10412 387852 10464
rect 72608 10344 72660 10396
rect 215484 10344 215536 10396
rect 240232 10344 240284 10396
rect 390652 10344 390704 10396
rect 69112 10276 69164 10328
rect 215392 10276 215444 10328
rect 255504 10276 255556 10328
rect 581736 10276 581788 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 156512 9392 156564 9444
rect 222568 9392 222620 9444
rect 234712 9392 234764 9444
rect 320916 9392 320968 9444
rect 149520 9324 149572 9376
rect 221280 9324 221332 9376
rect 236092 9324 236144 9376
rect 338672 9324 338724 9376
rect 142436 9256 142488 9308
rect 221188 9256 221240 9308
rect 236000 9256 236052 9308
rect 342168 9256 342220 9308
rect 62028 9188 62080 9240
rect 214196 9188 214248 9240
rect 237656 9188 237708 9240
rect 352840 9188 352892 9240
rect 54944 9120 54996 9172
rect 214104 9120 214156 9172
rect 237472 9120 237524 9172
rect 356336 9120 356388 9172
rect 7656 9052 7708 9104
rect 210792 9052 210844 9104
rect 237564 9052 237616 9104
rect 359924 9052 359976 9104
rect 2872 8984 2924 9036
rect 209964 8984 210016 9036
rect 261484 8984 261536 9036
rect 475752 8984 475804 9036
rect 1676 8916 1728 8968
rect 209872 8916 209924 8968
rect 254124 8916 254176 8968
rect 566832 8916 566884 8968
rect 202696 7964 202748 8016
rect 225236 7964 225288 8016
rect 195612 7896 195664 7948
rect 225328 7896 225380 7948
rect 167184 7828 167236 7880
rect 222476 7828 222528 7880
rect 230848 7828 230900 7880
rect 268844 7828 268896 7880
rect 158904 7760 158956 7812
rect 222384 7760 222436 7812
rect 232044 7760 232096 7812
rect 288992 7760 289044 7812
rect 148324 7692 148376 7744
rect 221004 7692 221056 7744
rect 233332 7692 233384 7744
rect 303160 7692 303212 7744
rect 144736 7624 144788 7676
rect 221096 7624 221148 7676
rect 257436 7624 257488 7676
rect 422576 7624 422628 7676
rect 121092 7556 121144 7608
rect 217324 7556 217376 7608
rect 257528 7556 257580 7608
rect 429660 7556 429712 7608
rect 230756 6672 230808 6724
rect 265348 6672 265400 6724
rect 187332 6604 187384 6656
rect 223764 6604 223816 6656
rect 230572 6604 230624 6656
rect 267740 6604 267792 6656
rect 183744 6536 183796 6588
rect 224408 6536 224460 6588
rect 230664 6536 230716 6588
rect 271236 6536 271288 6588
rect 180248 6468 180300 6520
rect 223856 6468 223908 6520
rect 231860 6468 231912 6520
rect 285404 6468 285456 6520
rect 176660 6400 176712 6452
rect 223948 6400 224000 6452
rect 241520 6400 241572 6452
rect 404820 6400 404872 6452
rect 130568 6332 130620 6384
rect 219808 6332 219860 6384
rect 241612 6332 241664 6384
rect 411904 6332 411956 6384
rect 117596 6264 117648 6316
rect 208032 6264 208084 6316
rect 231952 6264 232004 6316
rect 281908 6264 281960 6316
rect 282184 6264 282236 6316
rect 581000 6264 581052 6316
rect 92756 6196 92808 6248
rect 217508 6196 217560 6248
rect 253940 6196 253992 6248
rect 569132 6196 569184 6248
rect 25320 6128 25372 6180
rect 188344 6128 188396 6180
rect 197912 6128 197964 6180
rect 225144 6128 225196 6180
rect 254032 6128 254084 6180
rect 572720 6128 572772 6180
rect 201408 5380 201460 5432
rect 223488 5380 223540 5432
rect 187700 5312 187752 5364
rect 219624 5312 219676 5364
rect 162492 5244 162544 5296
rect 222936 5244 222988 5296
rect 150624 5176 150676 5228
rect 220912 5176 220964 5228
rect 147128 5108 147180 5160
rect 221556 5108 221608 5160
rect 237380 5108 237432 5160
rect 355232 5108 355284 5160
rect 127072 5040 127124 5092
rect 219716 5040 219768 5092
rect 248420 5040 248472 5092
rect 501788 5040 501840 5092
rect 110512 4972 110564 5024
rect 207940 4972 207992 5024
rect 251272 4972 251324 5024
rect 537208 4972 537260 5024
rect 60832 4904 60884 4956
rect 213920 4904 213972 4956
rect 230480 4904 230532 4956
rect 239404 4904 239456 4956
rect 252652 4904 252704 4956
rect 547880 4904 547932 4956
rect 15936 4836 15988 4888
rect 42064 4836 42116 4888
rect 58440 4836 58492 4888
rect 214012 4836 214064 4888
rect 214472 4836 214524 4888
rect 226616 4836 226668 4888
rect 229560 4836 229612 4888
rect 248788 4836 248840 4888
rect 252560 4836 252612 4888
rect 551468 4836 551520 4888
rect 32404 4768 32456 4820
rect 206284 4768 206336 4820
rect 210976 4768 211028 4820
rect 226524 4768 226576 4820
rect 229652 4768 229704 4820
rect 251180 4768 251232 4820
rect 255412 4768 255464 4820
rect 578608 4768 578660 4820
rect 200304 4088 200356 4140
rect 225696 4088 225748 4140
rect 185032 4020 185084 4072
rect 210424 4020 210476 4072
rect 219256 4020 219308 4072
rect 220820 4020 220872 4072
rect 177856 3952 177908 4004
rect 204904 3952 204956 4004
rect 233884 3952 233936 4004
rect 245200 3952 245252 4004
rect 132960 3884 133012 3936
rect 187700 3884 187752 3936
rect 193220 3884 193272 3936
rect 225052 3884 225104 3936
rect 229468 3884 229520 3936
rect 242900 3884 242952 3936
rect 104532 3816 104584 3868
rect 159364 3816 159416 3868
rect 166080 3816 166132 3868
rect 201408 3816 201460 3868
rect 218060 3816 218112 3868
rect 227352 3816 227404 3868
rect 229192 3816 229244 3868
rect 239220 3816 239272 3868
rect 239404 3816 239456 3868
rect 84476 3748 84528 3800
rect 140044 3748 140096 3800
rect 168472 3748 168524 3800
rect 213184 3748 213236 3800
rect 257620 3816 257672 3868
rect 264152 3816 264204 3868
rect 261760 3748 261812 3800
rect 276020 3748 276072 3800
rect 276756 3748 276808 3800
rect 106924 3680 106976 3732
rect 163504 3680 163556 3732
rect 179052 3680 179104 3732
rect 224224 3680 224276 3732
rect 228272 3680 228324 3732
rect 229836 3680 229888 3732
rect 99840 3612 99892 3664
rect 156604 3612 156656 3664
rect 161296 3612 161348 3664
rect 207664 3612 207716 3664
rect 216864 3612 216916 3664
rect 222292 3612 222344 3664
rect 227904 3612 227956 3664
rect 232228 3612 232280 3664
rect 233240 3612 233292 3664
rect 296076 3680 296128 3732
rect 307852 3680 307904 3732
rect 309048 3680 309100 3732
rect 316132 3680 316184 3732
rect 317328 3680 317380 3732
rect 236644 3612 236696 3664
rect 257068 3612 257120 3664
rect 257344 3612 257396 3664
rect 458088 3612 458140 3664
rect 93860 3544 93912 3596
rect 94780 3544 94832 3596
rect 102140 3544 102192 3596
rect 103336 3544 103388 3596
rect 110420 3544 110472 3596
rect 111616 3544 111668 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 125876 3544 125928 3596
rect 209044 3544 209096 3596
rect 209780 3544 209832 3596
rect 213276 3544 213328 3596
rect 229284 3544 229336 3596
rect 253480 3544 253532 3596
rect 255964 3544 256016 3596
rect 472256 3544 472308 3596
rect 473360 3544 473412 3596
rect 474188 3544 474240 3596
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 70308 3476 70360 3528
rect 30104 3408 30156 3460
rect 126980 3476 127032 3528
rect 128176 3476 128228 3528
rect 129372 3476 129424 3528
rect 219532 3476 219584 3528
rect 226340 3476 226392 3528
rect 228180 3476 228232 3528
rect 230112 3476 230164 3528
rect 244096 3476 244148 3528
rect 248052 3476 248104 3528
rect 484032 3544 484084 3596
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 127624 3408 127676 3460
rect 207756 3408 207808 3460
rect 229376 3408 229428 3460
rect 246396 3408 246448 3460
rect 252468 3408 252520 3460
rect 530124 3408 530176 3460
rect 168380 3340 168432 3392
rect 169576 3340 169628 3392
rect 184940 3340 184992 3392
rect 186136 3340 186188 3392
rect 190828 3340 190880 3392
rect 207848 3340 207900 3392
rect 227996 3340 228048 3392
rect 231032 3340 231084 3392
rect 231124 3340 231176 3392
rect 237012 3340 237064 3392
rect 239220 3340 239272 3392
rect 247592 3340 247644 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365812 3340 365864 3392
rect 367008 3340 367060 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 223948 3136 224000 3188
rect 228088 3136 228140 3188
rect 213368 3000 213420 3052
rect 220084 3000 220136 3052
rect 221556 3000 221608 3052
rect 227168 3000 227220 3052
rect 249984 3000 250036 3052
rect 256700 3000 256752 3052
rect 225144 2932 225196 2984
rect 226432 2932 226484 2984
rect 423680 1640 423732 1692
rect 424968 1640 425020 1692
rect 448520 1640 448572 1692
rect 449808 1640 449860 1692
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700398 40540 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 33784 700392 33836 700398
rect 33784 700334 33836 700340
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 51724 700392 51776 700398
rect 51724 700334 51776 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 15844 683188 15896 683194
rect 15844 683130 15896 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 4804 657008 4856 657014
rect 4804 656950 4856 656956
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3146 606112 3202 606121
rect 3146 606047 3202 606056
rect 3160 605946 3188 606047
rect 3148 605940 3200 605946
rect 3148 605882 3200 605888
rect 2778 580000 2834 580009
rect 2778 579935 2780 579944
rect 2832 579935 2834 579944
rect 2780 579906 2832 579912
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553586 3372 553823
rect 3332 553580 3384 553586
rect 3332 553522 3384 553528
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527270 2820 527847
rect 2780 527264 2832 527270
rect 2780 527206 2832 527212
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3436 466154 3464 619103
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 480254 3556 566879
rect 3528 480226 3648 480254
rect 3436 466126 3556 466154
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3436 462398 3464 462567
rect 3424 462392 3476 462398
rect 3424 462334 3476 462340
rect 3528 461786 3556 466126
rect 3516 461780 3568 461786
rect 3516 461722 3568 461728
rect 3620 457570 3648 480226
rect 3608 457564 3660 457570
rect 3608 457506 3660 457512
rect 4816 453354 4844 656950
rect 6184 605940 6236 605946
rect 6184 605882 6236 605888
rect 4896 579964 4948 579970
rect 4896 579906 4948 579912
rect 4804 453348 4856 453354
rect 4804 453290 4856 453296
rect 4908 450566 4936 579906
rect 4988 527264 5040 527270
rect 4988 527206 5040 527212
rect 5000 451926 5028 527206
rect 4988 451920 5040 451926
rect 4988 451862 5040 451868
rect 6196 450634 6224 605882
rect 7564 553580 7616 553586
rect 7564 553522 7616 553528
rect 7576 454714 7604 553522
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 14476 457638 14504 514762
rect 15856 475386 15884 683130
rect 15936 501016 15988 501022
rect 15936 500958 15988 500964
rect 15844 475380 15896 475386
rect 15844 475322 15896 475328
rect 14556 474768 14608 474774
rect 14556 474710 14608 474716
rect 14464 457632 14516 457638
rect 14464 457574 14516 457580
rect 7564 454708 7616 454714
rect 7564 454650 7616 454656
rect 14568 451994 14596 474710
rect 15948 454782 15976 500958
rect 15936 454776 15988 454782
rect 15936 454718 15988 454724
rect 14556 451988 14608 451994
rect 14556 451930 14608 451936
rect 6184 450628 6236 450634
rect 6184 450570 6236 450576
rect 4896 450560 4948 450566
rect 4896 450502 4948 450508
rect 2870 449576 2926 449585
rect 2870 449511 2926 449520
rect 2884 447846 2912 449511
rect 33796 448526 33824 700334
rect 37924 670744 37976 670750
rect 37924 670686 37976 670692
rect 37936 455394 37964 670686
rect 51736 463146 51764 700334
rect 55864 700324 55916 700330
rect 55864 700266 55916 700272
rect 51816 632120 51868 632126
rect 51816 632062 51868 632068
rect 51828 475454 51856 632062
rect 51816 475448 51868 475454
rect 51816 475390 51868 475396
rect 51724 463140 51776 463146
rect 51724 463082 51776 463088
rect 37924 455388 37976 455394
rect 37924 455330 37976 455336
rect 55876 452062 55904 700266
rect 71792 453422 71820 702986
rect 89180 700330 89208 703520
rect 105464 700398 105492 703520
rect 137848 700466 137876 703520
rect 154132 700534 154160 703520
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 170324 699718 170352 703520
rect 177396 700528 177448 700534
rect 177396 700470 177448 700476
rect 173256 700460 173308 700466
rect 173256 700402 173308 700408
rect 171784 700324 171836 700330
rect 171784 700266 171836 700272
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 78586 636440 78642 636449
rect 78586 636375 78642 636384
rect 78310 635352 78366 635361
rect 78310 635287 78366 635296
rect 78218 633720 78274 633729
rect 78218 633655 78274 633664
rect 77942 632632 77998 632641
rect 77942 632567 77998 632576
rect 77758 629640 77814 629649
rect 77758 629575 77814 629584
rect 77574 523288 77630 523297
rect 77574 523223 77630 523232
rect 77588 489598 77616 523223
rect 77772 520305 77800 629575
rect 77850 608696 77906 608705
rect 77850 608631 77906 608640
rect 77758 520296 77814 520305
rect 77758 520231 77814 520240
rect 77666 498400 77722 498409
rect 77666 498335 77722 498344
rect 77576 489592 77628 489598
rect 77576 489534 77628 489540
rect 77680 489462 77708 498335
rect 77772 489734 77800 520231
rect 77864 518894 77892 608631
rect 77956 523297 77984 632567
rect 78126 631000 78182 631009
rect 78126 630935 78182 630944
rect 78034 628008 78090 628017
rect 78034 627943 78090 627952
rect 78048 599962 78076 627943
rect 78140 600030 78168 630935
rect 78128 600024 78180 600030
rect 78128 599966 78180 599972
rect 78036 599956 78088 599962
rect 78036 599898 78088 599904
rect 78232 599894 78260 633655
rect 78220 599888 78272 599894
rect 78220 599830 78272 599836
rect 78324 584458 78352 635287
rect 78600 615494 78628 636375
rect 78508 615466 78628 615494
rect 78402 610056 78458 610065
rect 78402 609991 78458 610000
rect 78416 599758 78444 609991
rect 78404 599752 78456 599758
rect 78404 599694 78456 599700
rect 78508 599690 78536 615466
rect 78586 607744 78642 607753
rect 78586 607679 78642 607688
rect 78600 599826 78628 607679
rect 78588 599820 78640 599826
rect 78588 599762 78640 599768
rect 78496 599684 78548 599690
rect 78496 599626 78548 599632
rect 115848 597576 115900 597582
rect 103150 597544 103206 597553
rect 103150 597479 103206 597488
rect 111706 597544 111762 597553
rect 111706 597479 111762 597488
rect 115846 597544 115848 597553
rect 115900 597544 115902 597553
rect 115846 597479 115902 597488
rect 121366 597544 121422 597553
rect 121366 597479 121422 597488
rect 126886 597544 126942 597553
rect 126886 597479 126888 597488
rect 92478 597408 92534 597417
rect 92478 597343 92534 597352
rect 92492 596358 92520 597343
rect 103164 597310 103192 597479
rect 111720 597378 111748 597479
rect 111708 597372 111760 597378
rect 111708 597314 111760 597320
rect 103152 597304 103204 597310
rect 103152 597246 103204 597252
rect 94042 597136 94098 597145
rect 94042 597071 94098 597080
rect 103426 597136 103482 597145
rect 103426 597071 103482 597080
rect 106186 597136 106242 597145
rect 106186 597071 106188 597080
rect 79784 596352 79836 596358
rect 79784 596294 79836 596300
rect 92480 596352 92532 596358
rect 92480 596294 92532 596300
rect 78312 584452 78364 584458
rect 78312 584394 78364 584400
rect 78324 526561 78352 584394
rect 78494 526688 78550 526697
rect 78494 526623 78550 526632
rect 78310 526552 78366 526561
rect 78310 526487 78366 526496
rect 78310 523696 78366 523705
rect 78310 523631 78366 523640
rect 77942 523288 77998 523297
rect 77942 523223 77998 523232
rect 78126 520976 78182 520985
rect 78126 520911 78182 520920
rect 77864 518866 77984 518894
rect 77956 498681 77984 518866
rect 78034 517984 78090 517993
rect 78034 517919 78090 517928
rect 77942 498672 77998 498681
rect 77942 498607 77998 498616
rect 77760 489728 77812 489734
rect 77760 489670 77812 489676
rect 77668 489456 77720 489462
rect 77668 489398 77720 489404
rect 77956 467226 77984 498607
rect 78048 489802 78076 517919
rect 78140 489870 78168 520911
rect 78128 489864 78180 489870
rect 78128 489806 78180 489812
rect 78036 489796 78088 489802
rect 78036 489738 78088 489744
rect 78324 489666 78352 523631
rect 78312 489660 78364 489666
rect 78312 489602 78364 489608
rect 78508 489530 78536 526623
rect 78586 499896 78642 499905
rect 78586 499831 78642 499840
rect 78496 489524 78548 489530
rect 78496 489466 78548 489472
rect 78600 489394 78628 499831
rect 78588 489388 78640 489394
rect 78588 489330 78640 489336
rect 79796 488510 79824 596294
rect 94056 596290 94084 597071
rect 100666 597000 100722 597009
rect 100666 596935 100668 596944
rect 100720 596935 100722 596944
rect 100668 596906 100720 596912
rect 103440 596902 103468 597071
rect 106240 597071 106242 597080
rect 106188 597042 106240 597048
rect 121380 597038 121408 597479
rect 126940 597479 126942 597488
rect 131026 597544 131082 597553
rect 131026 597479 131082 597488
rect 136546 597544 136602 597553
rect 136546 597479 136602 597488
rect 140686 597544 140742 597553
rect 140686 597479 140742 597488
rect 126888 597450 126940 597456
rect 131040 597174 131068 597479
rect 136560 597446 136588 597479
rect 136548 597440 136600 597446
rect 136548 597382 136600 597388
rect 140700 597242 140728 597479
rect 140688 597236 140740 597242
rect 140688 597178 140740 597184
rect 131028 597168 131080 597174
rect 131028 597110 131080 597116
rect 121368 597032 121420 597038
rect 121368 596974 121420 596980
rect 103428 596896 103480 596902
rect 103428 596838 103480 596844
rect 104806 596864 104862 596873
rect 104806 596799 104808 596808
rect 104860 596799 104862 596808
rect 104808 596770 104860 596776
rect 95238 596320 95294 596329
rect 79876 596284 79928 596290
rect 79876 596226 79928 596232
rect 94044 596284 94096 596290
rect 95238 596255 95294 596264
rect 94044 596226 94096 596232
rect 79784 488504 79836 488510
rect 79784 488446 79836 488452
rect 79888 488442 79916 596226
rect 95252 596222 95280 596255
rect 79968 596216 80020 596222
rect 79968 596158 80020 596164
rect 95240 596216 95292 596222
rect 95240 596158 95292 596164
rect 79876 488436 79928 488442
rect 79876 488378 79928 488384
rect 79980 488374 80008 596158
rect 110510 489424 110566 489433
rect 110510 489359 110566 489368
rect 110524 488850 110552 489359
rect 110512 488844 110564 488850
rect 110512 488786 110564 488792
rect 120632 488708 120684 488714
rect 120632 488650 120684 488656
rect 115664 488640 115716 488646
rect 115664 488582 115716 488588
rect 105360 488572 105412 488578
rect 105360 488514 105412 488520
rect 92940 488504 92992 488510
rect 92938 488472 92940 488481
rect 105372 488481 105400 488514
rect 115676 488481 115704 488582
rect 120644 488481 120672 488650
rect 92992 488472 92994 488481
rect 92938 488407 92994 488416
rect 94226 488472 94282 488481
rect 94226 488407 94228 488416
rect 94280 488407 94282 488416
rect 97814 488472 97870 488481
rect 97814 488407 97870 488416
rect 99194 488472 99250 488481
rect 99194 488407 99250 488416
rect 100022 488472 100078 488481
rect 100022 488407 100078 488416
rect 101126 488472 101182 488481
rect 101126 488407 101182 488416
rect 102414 488472 102470 488481
rect 102414 488407 102470 488416
rect 104806 488472 104862 488481
rect 104806 488407 104862 488416
rect 105358 488472 105414 488481
rect 105358 488407 105414 488416
rect 105726 488472 105782 488481
rect 105726 488407 105782 488416
rect 115662 488472 115718 488481
rect 115662 488407 115718 488416
rect 120630 488472 120686 488481
rect 120630 488407 120686 488416
rect 125598 488472 125654 488481
rect 125598 488407 125654 488416
rect 130658 488472 130714 488481
rect 130658 488407 130714 488416
rect 135534 488472 135590 488481
rect 135534 488407 135590 488416
rect 140686 488472 140742 488481
rect 140686 488407 140742 488416
rect 94228 488378 94280 488384
rect 79968 488368 80020 488374
rect 95332 488368 95384 488374
rect 79968 488310 80020 488316
rect 95330 488336 95332 488345
rect 95384 488336 95386 488345
rect 95330 488271 95386 488280
rect 97828 487762 97856 488407
rect 97816 487756 97868 487762
rect 97816 487698 97868 487704
rect 99208 487558 99236 488407
rect 99196 487552 99248 487558
rect 99196 487494 99248 487500
rect 100036 487490 100064 488407
rect 100024 487484 100076 487490
rect 100024 487426 100076 487432
rect 101140 487354 101168 488407
rect 102428 487966 102456 488407
rect 102416 487960 102468 487966
rect 102416 487902 102468 487908
rect 104820 487626 104848 488407
rect 105740 487694 105768 488407
rect 125612 487830 125640 488407
rect 125600 487824 125652 487830
rect 125600 487766 125652 487772
rect 105728 487688 105780 487694
rect 105728 487630 105780 487636
rect 104808 487620 104860 487626
rect 104808 487562 104860 487568
rect 103426 487520 103482 487529
rect 103426 487455 103482 487464
rect 103440 487422 103468 487455
rect 103428 487416 103480 487422
rect 103428 487358 103480 487364
rect 101128 487348 101180 487354
rect 101128 487290 101180 487296
rect 130672 487218 130700 488407
rect 135548 487898 135576 488407
rect 135536 487892 135588 487898
rect 135536 487834 135588 487840
rect 140700 487286 140728 488407
rect 140688 487280 140740 487286
rect 140688 487222 140740 487228
rect 130660 487212 130712 487218
rect 130660 487154 130712 487160
rect 77944 467220 77996 467226
rect 77944 467162 77996 467168
rect 71780 453416 71832 453422
rect 71780 453358 71832 453364
rect 55864 452056 55916 452062
rect 55864 451998 55916 452004
rect 33784 448520 33836 448526
rect 33784 448462 33836 448468
rect 171796 447914 171824 700266
rect 173164 699712 173216 699718
rect 173164 699654 173216 699660
rect 173176 450770 173204 699654
rect 173268 475522 173296 700402
rect 177304 700392 177356 700398
rect 177304 700334 177356 700340
rect 173256 475516 173308 475522
rect 173256 475458 173308 475464
rect 177316 452130 177344 700334
rect 177408 471306 177436 700470
rect 202800 700466 202828 703520
rect 188988 700460 189040 700466
rect 188988 700402 189040 700408
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 186870 637120 186926 637129
rect 186870 637055 186926 637064
rect 186778 636032 186834 636041
rect 186778 635967 186834 635976
rect 186594 608424 186650 608433
rect 186594 608359 186650 608368
rect 186608 599826 186636 608359
rect 186596 599820 186648 599826
rect 186596 599762 186648 599768
rect 186608 498273 186636 599762
rect 186792 586514 186820 635967
rect 186884 599690 186912 637055
rect 187330 634400 187386 634409
rect 187330 634335 187386 634344
rect 187238 631680 187294 631689
rect 187238 631615 187294 631624
rect 187146 628688 187202 628697
rect 187146 628623 187202 628632
rect 187054 610328 187110 610337
rect 187054 610263 187110 610272
rect 187068 599758 187096 610263
rect 187160 599962 187188 628623
rect 187252 600030 187280 631615
rect 187240 600024 187292 600030
rect 187240 599966 187292 599972
rect 187148 599956 187200 599962
rect 187148 599898 187200 599904
rect 187056 599752 187108 599758
rect 187056 599694 187108 599700
rect 186872 599684 186924 599690
rect 186872 599626 186924 599632
rect 186700 586486 186820 586514
rect 186700 584458 186728 586486
rect 186688 584452 186740 584458
rect 186688 584394 186740 584400
rect 186700 526017 186728 584394
rect 186884 527105 186912 599626
rect 186870 527096 186926 527105
rect 186870 527031 186926 527040
rect 186686 526008 186742 526017
rect 186686 525943 186742 525952
rect 186884 525910 186912 527031
rect 186872 525904 186924 525910
rect 186872 525846 186924 525852
rect 187068 500313 187096 599694
rect 187160 518430 187188 599898
rect 187252 521665 187280 599966
rect 187344 599894 187372 634335
rect 187422 633312 187478 633321
rect 187422 633247 187478 633256
rect 187332 599888 187384 599894
rect 187332 599830 187384 599836
rect 187344 524385 187372 599830
rect 187330 524376 187386 524385
rect 187330 524311 187386 524320
rect 187436 523297 187464 633247
rect 187514 630320 187570 630329
rect 187514 630255 187570 630264
rect 187422 523288 187478 523297
rect 187422 523223 187478 523232
rect 187238 521656 187294 521665
rect 187528 521626 187556 630255
rect 187606 608696 187662 608705
rect 187606 608631 187662 608640
rect 187238 521591 187294 521600
rect 187516 521620 187568 521626
rect 187516 521562 187568 521568
rect 187148 518424 187200 518430
rect 187148 518366 187200 518372
rect 187054 500304 187110 500313
rect 187054 500239 187110 500248
rect 187068 499574 187096 500239
rect 186976 499546 187096 499574
rect 186594 498264 186650 498273
rect 186594 498199 186650 498208
rect 186976 489394 187004 499546
rect 187620 498681 187648 608631
rect 188712 596352 188764 596358
rect 188712 596294 188764 596300
rect 187700 525904 187752 525910
rect 187700 525846 187752 525852
rect 187606 498672 187662 498681
rect 187606 498607 187662 498616
rect 187054 498264 187110 498273
rect 187054 498199 187110 498208
rect 187068 489462 187096 498199
rect 187056 489456 187108 489462
rect 187056 489398 187108 489404
rect 186964 489388 187016 489394
rect 186964 489330 187016 489336
rect 177396 471300 177448 471306
rect 177396 471242 177448 471248
rect 186976 469198 187004 489330
rect 187068 485110 187096 489398
rect 187056 485104 187108 485110
rect 187056 485046 187108 485052
rect 187620 476814 187648 498607
rect 187712 489530 187740 525846
rect 188342 524376 188398 524385
rect 188342 524311 188398 524320
rect 187790 523288 187846 523297
rect 187790 523223 187846 523232
rect 187804 489598 187832 523223
rect 187974 521656 188030 521665
rect 187974 521591 188030 521600
rect 188160 521620 188212 521626
rect 187988 489870 188016 521591
rect 188160 521562 188212 521568
rect 188172 520305 188200 521562
rect 188158 520296 188214 520305
rect 188158 520231 188214 520240
rect 188066 518664 188122 518673
rect 188066 518599 188122 518608
rect 188080 518430 188108 518599
rect 188068 518424 188120 518430
rect 188068 518366 188120 518372
rect 187976 489864 188028 489870
rect 187976 489806 188028 489812
rect 187792 489592 187844 489598
rect 187792 489534 187844 489540
rect 187700 489524 187752 489530
rect 187700 489466 187752 489472
rect 187712 486470 187740 489466
rect 187804 488782 187832 489534
rect 187988 488918 188016 489806
rect 188080 489802 188108 518366
rect 188068 489796 188120 489802
rect 188068 489738 188120 489744
rect 187976 488912 188028 488918
rect 187976 488854 188028 488860
rect 188080 488866 188108 489738
rect 188172 489734 188200 520231
rect 188160 489728 188212 489734
rect 188160 489670 188212 489676
rect 188172 489002 188200 489670
rect 188356 489666 188384 524311
rect 188344 489660 188396 489666
rect 188344 489602 188396 489608
rect 188356 489190 188384 489602
rect 188344 489184 188396 489190
rect 188344 489126 188396 489132
rect 188172 488974 188568 489002
rect 188080 488838 188384 488866
rect 187792 488776 187844 488782
rect 187792 488718 187844 488724
rect 188252 488776 188304 488782
rect 188252 488718 188304 488724
rect 187700 486464 187752 486470
rect 187700 486406 187752 486412
rect 188264 478174 188292 488718
rect 188252 478168 188304 478174
rect 188252 478110 188304 478116
rect 187608 476808 187660 476814
rect 187608 476750 187660 476756
rect 188356 473346 188384 488838
rect 188540 474706 188568 488974
rect 188620 488912 188672 488918
rect 188620 488854 188672 488860
rect 188632 477494 188660 488854
rect 188724 488510 188752 596294
rect 188896 596284 188948 596290
rect 188896 596226 188948 596232
rect 188804 596216 188856 596222
rect 188804 596158 188856 596164
rect 188712 488504 188764 488510
rect 188712 488446 188764 488452
rect 188724 488102 188752 488446
rect 188816 488442 188844 596158
rect 188804 488436 188856 488442
rect 188804 488378 188856 488384
rect 188712 488096 188764 488102
rect 188712 488038 188764 488044
rect 188816 488034 188844 488378
rect 188908 488345 188936 596226
rect 188894 488336 188950 488345
rect 188894 488271 188950 488280
rect 188804 488028 188856 488034
rect 188804 487970 188856 487976
rect 188620 477488 188672 477494
rect 188620 477430 188672 477436
rect 188528 474700 188580 474706
rect 188528 474642 188580 474648
rect 188344 473340 188396 473346
rect 188344 473282 188396 473288
rect 186964 469192 187016 469198
rect 186964 469134 187016 469140
rect 177304 452124 177356 452130
rect 177304 452066 177356 452072
rect 173164 450764 173216 450770
rect 173164 450706 173216 450712
rect 171784 447908 171836 447914
rect 171784 447850 171836 447856
rect 2872 447840 2924 447846
rect 2872 447782 2924 447788
rect 6184 446548 6236 446554
rect 6184 446490 6236 446496
rect 3700 445052 3752 445058
rect 3700 444994 3752 445000
rect 3608 443692 3660 443698
rect 3608 443634 3660 443640
rect 3424 443012 3476 443018
rect 3424 442954 3476 442960
rect 3056 372564 3108 372570
rect 3056 372506 3108 372512
rect 3068 371385 3096 372506
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 2780 320136 2832 320142
rect 2780 320078 2832 320084
rect 2792 319297 2820 320078
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3240 293956 3292 293962
rect 3240 293898 3292 293904
rect 3252 293185 3280 293898
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3148 254788 3200 254794
rect 3148 254730 3200 254736
rect 3160 254153 3188 254730
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3332 241460 3384 241466
rect 3332 241402 3384 241408
rect 3344 241097 3372 241402
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3148 215280 3200 215286
rect 3148 215222 3200 215228
rect 3160 214985 3188 215222
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3332 59356 3384 59362
rect 3332 59298 3384 59304
rect 3344 58585 3372 59298
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3436 45529 3464 442954
rect 3516 423632 3568 423638
rect 3514 423600 3516 423609
rect 3568 423600 3570 423609
rect 3514 423535 3570 423544
rect 3516 411256 3568 411262
rect 3516 411198 3568 411204
rect 3528 410553 3556 411198
rect 3514 410544 3570 410553
rect 3514 410479 3570 410488
rect 3516 398812 3568 398818
rect 3516 398754 3568 398760
rect 3528 397497 3556 398754
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3516 358760 3568 358766
rect 3516 358702 3568 358708
rect 3528 358465 3556 358702
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3516 352572 3568 352578
rect 3516 352514 3568 352520
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3436 32473 3464 32982
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 13116 3476 13122
rect 3424 13058 3476 13064
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 570 4856 626 4865
rect 570 4791 626 4800
rect 584 480 612 4791
rect 1688 480 1716 8910
rect 2884 480 2912 8978
rect 3436 490 3464 13058
rect 3528 6497 3556 352514
rect 3620 136785 3648 443634
rect 3712 188873 3740 444994
rect 4160 351212 4212 351218
rect 4160 351154 4212 351160
rect 3698 188864 3754 188873
rect 3698 188799 3754 188808
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 4172 16574 4200 351154
rect 6196 254794 6224 446490
rect 189000 446486 189028 700402
rect 218992 700398 219020 703520
rect 190000 700392 190052 700398
rect 190000 700334 190052 700340
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 189908 700324 189960 700330
rect 189908 700266 189960 700272
rect 189078 526008 189134 526017
rect 189078 525943 189134 525952
rect 189092 478854 189120 525943
rect 189920 487801 189948 700266
rect 189906 487792 189962 487801
rect 189906 487727 189962 487736
rect 189080 478848 189132 478854
rect 189080 478790 189132 478796
rect 188988 446480 189040 446486
rect 188988 446422 189040 446428
rect 190012 446418 190040 700334
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 281540 700324 281592 700330
rect 281540 700266 281592 700272
rect 225512 597576 225564 597582
rect 209962 597544 210018 597553
rect 209962 597479 210018 597488
rect 212354 597544 212410 597553
rect 212354 597479 212410 597488
rect 213826 597544 213882 597553
rect 213826 597479 213882 597488
rect 214838 597544 214894 597553
rect 214838 597479 214894 597488
rect 215298 597544 215354 597553
rect 215298 597479 215354 597488
rect 219438 597544 219494 597553
rect 219438 597479 219494 597488
rect 225510 597544 225512 597553
rect 225564 597544 225566 597553
rect 225510 597479 225566 597488
rect 230662 597544 230718 597553
rect 230662 597479 230718 597488
rect 234618 597544 234674 597553
rect 234618 597479 234620 597488
rect 209042 597408 209098 597417
rect 209042 597343 209098 597352
rect 207662 597272 207718 597281
rect 207662 597207 207718 597216
rect 204350 596592 204406 596601
rect 204350 596527 204406 596536
rect 202878 596456 202934 596465
rect 202878 596391 202934 596400
rect 202892 596358 202920 596391
rect 202880 596352 202932 596358
rect 202880 596294 202932 596300
rect 204258 596320 204314 596329
rect 204364 596290 204392 596527
rect 207676 596290 207704 597207
rect 209056 596358 209084 597343
rect 209976 596970 210004 597479
rect 212368 597310 212396 597479
rect 212356 597304 212408 597310
rect 212356 597246 212408 597252
rect 209964 596964 210016 596970
rect 209964 596906 210016 596912
rect 211068 596964 211120 596970
rect 211068 596906 211120 596912
rect 211080 596426 211108 596906
rect 211068 596420 211120 596426
rect 211068 596362 211120 596368
rect 209044 596352 209096 596358
rect 209044 596294 209096 596300
rect 204258 596255 204314 596264
rect 204352 596284 204404 596290
rect 204272 596222 204300 596255
rect 204352 596226 204404 596232
rect 207664 596284 207716 596290
rect 207664 596226 207716 596232
rect 212368 596222 212396 597246
rect 212446 597000 212502 597009
rect 212446 596935 212502 596944
rect 212460 596494 212488 596935
rect 213840 596902 213868 597479
rect 213828 596896 213880 596902
rect 213828 596838 213880 596844
rect 213840 596562 213868 596838
rect 214852 596834 214880 597479
rect 215312 597106 215340 597479
rect 219452 597378 219480 597479
rect 219440 597372 219492 597378
rect 219440 597314 219492 597320
rect 220728 597372 220780 597378
rect 220728 597314 220780 597320
rect 215300 597100 215352 597106
rect 215300 597042 215352 597048
rect 214840 596828 214892 596834
rect 214840 596770 214892 596776
rect 214852 596630 214880 596770
rect 215312 596698 215340 597042
rect 220740 596766 220768 597314
rect 230676 596834 230704 597479
rect 234672 597479 234674 597488
rect 240506 597544 240562 597553
rect 240506 597479 240562 597488
rect 245474 597544 245530 597553
rect 245474 597479 245530 597488
rect 250534 597544 250590 597553
rect 250534 597479 250590 597488
rect 234620 597450 234672 597456
rect 234632 596902 234660 597450
rect 240520 596970 240548 597479
rect 245488 597446 245516 597479
rect 245476 597440 245528 597446
rect 245476 597382 245528 597388
rect 250548 597106 250576 597479
rect 250536 597100 250588 597106
rect 250536 597042 250588 597048
rect 240508 596964 240560 596970
rect 240508 596906 240560 596912
rect 234620 596896 234672 596902
rect 234620 596838 234672 596844
rect 230664 596828 230716 596834
rect 230664 596770 230716 596776
rect 220728 596760 220780 596766
rect 220728 596702 220780 596708
rect 280988 596760 281040 596766
rect 280988 596702 281040 596708
rect 215300 596692 215352 596698
rect 215300 596634 215352 596640
rect 214840 596624 214892 596630
rect 214840 596566 214892 596572
rect 213828 596556 213880 596562
rect 213828 596498 213880 596504
rect 212448 596488 212500 596494
rect 212448 596430 212500 596436
rect 204260 596216 204312 596222
rect 204260 596158 204312 596164
rect 212356 596216 212408 596222
rect 212356 596158 212408 596164
rect 240784 489184 240836 489190
rect 240784 489126 240836 489132
rect 220728 488844 220780 488850
rect 220728 488786 220780 488792
rect 215300 488776 215352 488782
rect 215300 488718 215352 488724
rect 215312 488578 215340 488718
rect 220740 488578 220768 488786
rect 230480 488708 230532 488714
rect 230480 488650 230532 488656
rect 231768 488708 231820 488714
rect 231768 488650 231820 488656
rect 226248 488640 226300 488646
rect 226248 488582 226300 488588
rect 215300 488572 215352 488578
rect 215300 488514 215352 488520
rect 220728 488572 220780 488578
rect 220728 488514 220780 488520
rect 215312 488481 215340 488514
rect 220740 488481 220768 488514
rect 226260 488481 226288 488582
rect 230492 488481 230520 488650
rect 231780 488510 231808 488650
rect 231768 488504 231820 488510
rect 215298 488472 215354 488481
rect 215298 488407 215354 488416
rect 220726 488472 220782 488481
rect 220726 488407 220782 488416
rect 226246 488472 226302 488481
rect 226246 488407 226302 488416
rect 230478 488472 230534 488481
rect 231768 488446 231820 488452
rect 230478 488407 230534 488416
rect 202880 488096 202932 488102
rect 202878 488064 202880 488073
rect 202932 488064 202934 488073
rect 202878 487999 202934 488008
rect 204258 488064 204314 488073
rect 204258 487999 204260 488008
rect 204312 487999 204314 488008
rect 211802 488064 211858 488073
rect 211802 487999 211858 488008
rect 204260 487970 204312 487976
rect 211816 487966 211844 487999
rect 211804 487960 211856 487966
rect 211158 487928 211214 487937
rect 211804 487902 211856 487908
rect 219624 487960 219676 487966
rect 219624 487902 219676 487908
rect 211158 487863 211214 487872
rect 207664 487756 207716 487762
rect 207664 487698 207716 487704
rect 204902 487384 204958 487393
rect 204902 487319 204958 487328
rect 203522 487248 203578 487257
rect 203522 487183 203578 487192
rect 203536 448458 203564 487183
rect 204916 459474 204944 487319
rect 207676 487257 207704 487698
rect 209044 487552 209096 487558
rect 209044 487494 209096 487500
rect 210054 487520 210110 487529
rect 209056 487257 209084 487494
rect 210054 487455 210056 487464
rect 210108 487455 210110 487464
rect 211068 487484 211120 487490
rect 210056 487426 210108 487432
rect 211068 487426 211120 487432
rect 205086 487248 205142 487257
rect 205086 487183 205142 487192
rect 207662 487248 207718 487257
rect 207662 487183 207718 487192
rect 209042 487248 209098 487257
rect 209042 487183 209098 487192
rect 204904 459468 204956 459474
rect 204904 459410 204956 459416
rect 205100 459406 205128 487183
rect 207676 481098 207704 487183
rect 207664 481092 207716 481098
rect 207664 481034 207716 481040
rect 205088 459400 205140 459406
rect 205088 459342 205140 459348
rect 209056 449818 209084 487183
rect 211080 482322 211108 487426
rect 211172 487354 211200 487863
rect 211160 487348 211212 487354
rect 211160 487290 211212 487296
rect 211160 484424 211212 484430
rect 211160 484366 211212 484372
rect 211068 482316 211120 482322
rect 211068 482258 211120 482264
rect 209044 449812 209096 449818
rect 209044 449754 209096 449760
rect 203524 448452 203576 448458
rect 203524 448394 203576 448400
rect 211172 446758 211200 484366
rect 211344 456816 211396 456822
rect 211344 456758 211396 456764
rect 211160 446752 211212 446758
rect 209594 446720 209650 446729
rect 204904 446684 204956 446690
rect 211160 446694 211212 446700
rect 209594 446655 209650 446664
rect 204904 446626 204956 446632
rect 190000 446412 190052 446418
rect 190000 446354 190052 446360
rect 200856 446344 200908 446350
rect 200856 446286 200908 446292
rect 204350 446312 204406 446321
rect 184204 446208 184256 446214
rect 184204 446150 184256 446156
rect 14464 445868 14516 445874
rect 14464 445810 14516 445816
rect 6276 445460 6328 445466
rect 6276 445402 6328 445408
rect 6288 320142 6316 445402
rect 11058 395312 11114 395321
rect 11058 395247 11114 395256
rect 6276 320136 6328 320142
rect 6276 320078 6328 320084
rect 6184 254788 6236 254794
rect 6184 254730 6236 254736
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5552 16574 5580 22714
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3436 462 3648 490
rect 5276 480 5304 16546
rect 3620 354 3648 462
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7668 480 7696 9046
rect 8772 480 8800 13126
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 15846
rect 11072 6914 11100 395247
rect 13820 354000 13872 354006
rect 11150 353968 11206 353977
rect 13820 353942 13872 353948
rect 11150 353903 11206 353912
rect 11164 16574 11192 353903
rect 13832 16574 13860 353942
rect 14476 306338 14504 445810
rect 106924 445392 106976 445398
rect 106924 445334 106976 445340
rect 35164 443080 35216 443086
rect 35164 443022 35216 443028
rect 35176 398818 35204 443022
rect 35164 398812 35216 398818
rect 35164 398754 35216 398760
rect 15844 398132 15896 398138
rect 15844 398074 15896 398080
rect 14464 306332 14516 306338
rect 14464 306274 14516 306280
rect 15856 22778 15884 398074
rect 42062 398032 42118 398041
rect 42062 397967 42118 397976
rect 37280 397316 37332 397322
rect 37280 397258 37332 397264
rect 27618 395448 27674 395457
rect 27618 395383 27674 395392
rect 23480 358080 23532 358086
rect 23480 358022 23532 358028
rect 19340 354136 19392 354142
rect 19340 354078 19392 354084
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 11164 16546 11928 16574
rect 13832 16546 14320 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13542 13016 13598 13025
rect 13542 12951 13598 12960
rect 13556 480 13584 12951
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17038 11656 17094 11665
rect 17038 11591 17094 11600
rect 15936 4888 15988 4894
rect 15936 4830 15988 4836
rect 15948 480 15976 4830
rect 17052 480 17080 11591
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 14418
rect 19352 3534 19380 354078
rect 19432 354068 19484 354074
rect 19432 354010 19484 354016
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19444 480 19472 354010
rect 23492 16574 23520 358022
rect 23492 16546 24256 16574
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20272 354 20300 3470
rect 21836 480 21864 11698
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 14486
rect 24228 480 24256 16546
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 25320 6180 25372 6186
rect 25320 6122 25372 6128
rect 25332 480 25360 6122
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 11766
rect 27632 3534 27660 395383
rect 34520 392624 34572 392630
rect 34520 392566 34572 392572
rect 30378 355328 30434 355337
rect 30378 355263 30434 355272
rect 30392 16574 30420 355263
rect 30392 16546 30880 16574
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 14554
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 30116 480 30144 3402
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 32416 480 32444 4762
rect 33612 480 33640 11834
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 392566
rect 37292 16574 37320 397258
rect 40040 396840 40092 396846
rect 40040 396782 40092 396788
rect 38660 175976 38712 175982
rect 38660 175918 38712 175924
rect 38672 16574 38700 175918
rect 40052 16574 40080 396782
rect 41420 354204 41472 354210
rect 41420 354146 41472 354152
rect 41432 16574 41460 354146
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35992 15972 36044 15978
rect 35992 15914 36044 15920
rect 36004 480 36032 15914
rect 36728 11960 36780 11966
rect 36728 11902 36780 11908
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 11902
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 42076 4894 42104 397967
rect 48318 396672 48374 396681
rect 48318 396607 48374 396616
rect 46938 393952 46994 393961
rect 46938 393887 46994 393896
rect 45560 355360 45612 355366
rect 45560 355302 45612 355308
rect 42800 354272 42852 354278
rect 42800 354214 42852 354220
rect 42064 4888 42116 4894
rect 42064 4830 42116 4836
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 354214
rect 45572 16574 45600 355302
rect 46952 16574 46980 393887
rect 48332 16574 48360 396607
rect 67638 395584 67694 395593
rect 67638 395519 67694 395528
rect 63500 393984 63552 393990
rect 63500 393926 63552 393932
rect 56600 354340 56652 354346
rect 56600 354282 56652 354288
rect 52460 352640 52512 352646
rect 52460 352582 52512 352588
rect 49698 351112 49754 351121
rect 49698 351047 49754 351056
rect 49712 16574 49740 351047
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44180 14680 44232 14686
rect 44180 14622 44232 14628
rect 44192 3534 44220 14622
rect 44272 12028 44324 12034
rect 44272 11970 44324 11976
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 11970
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51354 8936 51410 8945
rect 51354 8871 51410 8880
rect 51368 480 51396 8871
rect 52472 3534 52500 352582
rect 56612 16574 56640 354282
rect 63512 16574 63540 393926
rect 56612 16546 56824 16574
rect 63512 16546 64368 16574
rect 56048 13320 56100 13326
rect 56048 13262 56100 13268
rect 52552 13252 52604 13258
rect 52552 13194 52604 13200
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 13194
rect 54944 9172 54996 9178
rect 54944 9114 54996 9120
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 9114
rect 56060 480 56088 13262
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 63224 13456 63276 13462
rect 63224 13398 63276 13404
rect 59360 13388 59412 13394
rect 59360 13330 59412 13336
rect 58440 4888 58492 4894
rect 58440 4830 58492 4836
rect 58452 480 58480 4830
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13330
rect 62028 9240 62080 9246
rect 62028 9182 62080 9188
rect 60832 4956 60884 4962
rect 60832 4898 60884 4904
rect 60844 480 60872 4898
rect 62040 480 62068 9182
rect 63236 480 63264 13398
rect 64340 480 64368 16546
rect 66718 13152 66774 13161
rect 66718 13087 66774 13096
rect 65062 10296 65118 10305
rect 65062 10231 65118 10240
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 10231
rect 66732 480 66760 13087
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 395519
rect 93860 395480 93912 395486
rect 93860 395422 93912 395428
rect 86960 395412 87012 395418
rect 86960 395354 87012 395360
rect 77300 395344 77352 395350
rect 77300 395286 77352 395292
rect 73160 355428 73212 355434
rect 73160 355370 73212 355376
rect 73172 16574 73200 355370
rect 73172 16546 73384 16574
rect 71504 16040 71556 16046
rect 71504 15982 71556 15988
rect 69112 10328 69164 10334
rect 69112 10270 69164 10276
rect 69124 480 69152 10270
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 70320 480 70348 3470
rect 71516 480 71544 15982
rect 72608 10396 72660 10402
rect 72608 10338 72660 10344
rect 72620 480 72648 10338
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75000 14748 75052 14754
rect 75000 14690 75052 14696
rect 75012 480 75040 14690
rect 75920 10464 75972 10470
rect 75920 10406 75972 10412
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 10406
rect 77312 6914 77340 395286
rect 82818 394088 82874 394097
rect 82818 394023 82874 394032
rect 78680 354408 78732 354414
rect 78680 354350 78732 354356
rect 77392 177336 77444 177342
rect 77392 177278 77444 177284
rect 77404 16574 77432 177278
rect 78692 16574 78720 354350
rect 81438 177304 81494 177313
rect 81438 177239 81494 177248
rect 81452 16574 81480 177239
rect 82832 16574 82860 394023
rect 85578 177440 85634 177449
rect 85578 177375 85634 177384
rect 85592 16574 85620 177375
rect 86972 16574 87000 395354
rect 88340 355496 88392 355502
rect 88340 355438 88392 355444
rect 88352 16574 88380 355438
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80888 13524 80940 13530
rect 80888 13466 80940 13472
rect 80900 480 80928 13466
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84476 3800 84528 3806
rect 84476 3742 84528 3748
rect 84488 480 84516 3742
rect 85684 480 85712 16546
rect 86408 10532 86460 10538
rect 86408 10474 86460 10480
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 10474
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 91560 14816 91612 14822
rect 91560 14758 91612 14764
rect 89904 10600 89956 10606
rect 89904 10542 89956 10548
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 10542
rect 91572 480 91600 14758
rect 92756 6248 92808 6254
rect 92756 6190 92808 6196
rect 92768 480 92796 6190
rect 93872 3602 93900 395422
rect 106936 372570 106964 445334
rect 157984 444916 158036 444922
rect 157984 444858 158036 444864
rect 157996 423638 158024 444858
rect 157984 423632 158036 423638
rect 157984 423574 158036 423580
rect 171140 398268 171192 398274
rect 171140 398210 171192 398216
rect 139400 398200 139452 398206
rect 139400 398142 139452 398148
rect 131120 396908 131172 396914
rect 131120 396850 131172 396856
rect 121458 395856 121514 395865
rect 121458 395791 121514 395800
rect 118698 395720 118754 395729
rect 118698 395655 118754 395664
rect 115940 395616 115992 395622
rect 115940 395558 115992 395564
rect 109040 395548 109092 395554
rect 109040 395490 109092 395496
rect 106924 372564 106976 372570
rect 106924 372506 106976 372512
rect 104900 352708 104952 352714
rect 104900 352650 104952 352656
rect 102140 171828 102192 171834
rect 102140 171770 102192 171776
rect 95240 35216 95292 35222
rect 95240 35158 95292 35164
rect 95252 16574 95280 35158
rect 95252 16546 95832 16574
rect 93952 10668 94004 10674
rect 93952 10610 94004 10616
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93964 480 93992 10610
rect 94780 3596 94832 3602
rect 94780 3538 94832 3544
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94792 354 94820 3538
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 98184 14884 98236 14890
rect 98184 14826 98236 14832
rect 97448 10736 97500 10742
rect 97448 10678 97500 10684
rect 97460 480 97488 10678
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 14826
rect 100758 10432 100814 10441
rect 100758 10367 100814 10376
rect 99840 3664 99892 3670
rect 99840 3606 99892 3612
rect 99852 480 99880 3606
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 10367
rect 102152 3602 102180 171770
rect 104912 16574 104940 352650
rect 104912 16546 105768 16574
rect 102230 14512 102286 14521
rect 102230 14447 102286 14456
rect 102140 3596 102192 3602
rect 102140 3538 102192 3544
rect 102244 480 102272 14447
rect 104532 3868 104584 3874
rect 104532 3810 104584 3816
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 104544 480 104572 3810
rect 105740 480 105768 16546
rect 108120 12096 108172 12102
rect 108120 12038 108172 12044
rect 106924 3732 106976 3738
rect 106924 3674 106976 3680
rect 106936 480 106964 3674
rect 108132 480 108160 12038
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 395490
rect 113180 355564 113232 355570
rect 113180 355506 113232 355512
rect 113192 16574 113220 355506
rect 115952 16574 115980 395558
rect 113192 16546 114048 16574
rect 115952 16546 116440 16574
rect 112352 14952 112404 14958
rect 112352 14894 112404 14900
rect 110420 12164 110472 12170
rect 110420 12106 110472 12112
rect 110432 3602 110460 12106
rect 110512 5024 110564 5030
rect 110512 4966 110564 4972
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 110524 480 110552 4966
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111628 480 111656 3538
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 14894
rect 114020 480 114048 16546
rect 114744 12232 114796 12238
rect 114744 12174 114796 12180
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 12174
rect 116412 480 116440 16546
rect 117596 6316 117648 6322
rect 117596 6258 117648 6264
rect 117608 480 117636 6258
rect 118712 3602 118740 395655
rect 118790 351248 118846 351257
rect 118790 351183 118846 351192
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 118804 480 118832 351183
rect 121472 16574 121500 395791
rect 127622 354104 127678 354113
rect 127622 354039 127678 354048
rect 122838 352608 122894 352617
rect 122838 352543 122894 352552
rect 122852 16574 122880 352543
rect 126980 177404 127032 177410
rect 126980 177346 127032 177352
rect 124220 37936 124272 37942
rect 124220 37878 124272 37884
rect 124232 16574 124260 37878
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 121092 7608 121144 7614
rect 121092 7550 121144 7556
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 119908 480 119936 3538
rect 121104 480 121132 7550
rect 122300 480 122328 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 125888 480 125916 3538
rect 126992 3534 127020 177346
rect 127072 5092 127124 5098
rect 127072 5034 127124 5040
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 127084 2530 127112 5034
rect 127636 3466 127664 354039
rect 131132 16574 131160 396850
rect 138018 396808 138074 396817
rect 138018 396743 138074 396752
rect 135258 352744 135314 352753
rect 135258 352679 135314 352688
rect 133880 177472 133932 177478
rect 133880 177414 133932 177420
rect 131132 16546 131344 16574
rect 130568 6384 130620 6390
rect 130568 6326 130620 6332
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 127624 3460 127676 3466
rect 127624 3402 127676 3408
rect 126992 2502 127112 2530
rect 126992 480 127020 2502
rect 128188 480 128216 3470
rect 129384 480 129412 3470
rect 130580 480 130608 6326
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132960 3936 133012 3942
rect 132960 3878 133012 3884
rect 132972 480 133000 3878
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 177414
rect 135272 480 135300 352679
rect 138032 16574 138060 396743
rect 139412 16574 139440 398142
rect 162860 397112 162912 397118
rect 162860 397054 162912 397060
rect 151820 397044 151872 397050
rect 151820 396986 151872 396992
rect 144920 396976 144972 396982
rect 144920 396918 144972 396924
rect 143540 394052 143592 394058
rect 143540 393994 143592 394000
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 136456 16108 136508 16114
rect 136456 16050 136508 16056
rect 136468 480 136496 16050
rect 137650 7576 137706 7585
rect 137650 7511 137706 7520
rect 137664 480 137692 7511
rect 138860 480 138888 16546
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 140042 13288 140098 13297
rect 140042 13223 140098 13232
rect 140056 3806 140084 13223
rect 142436 9308 142488 9314
rect 142436 9250 142488 9256
rect 141238 7712 141294 7721
rect 141238 7647 141294 7656
rect 140044 3800 140096 3806
rect 140044 3742 140096 3748
rect 141252 480 141280 7647
rect 142448 480 142476 9250
rect 143552 480 143580 393994
rect 144932 16574 144960 396918
rect 144932 16546 145512 16574
rect 144736 7676 144788 7682
rect 144736 7618 144788 7624
rect 144748 480 144776 7618
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 151832 9674 151860 396986
rect 154578 394224 154634 394233
rect 154578 394159 154634 394168
rect 153198 351384 153254 351393
rect 153198 351319 153254 351328
rect 151912 351280 151964 351286
rect 151912 351222 151964 351228
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 149520 9376 149572 9382
rect 149520 9318 149572 9324
rect 148324 7744 148376 7750
rect 148324 7686 148376 7692
rect 147128 5160 147180 5166
rect 147128 5102 147180 5108
rect 147140 480 147168 5102
rect 148336 480 148364 7686
rect 149532 480 149560 9318
rect 151924 6914 151952 351222
rect 153212 16574 153240 351319
rect 154592 16574 154620 394159
rect 156602 354240 156658 354249
rect 156602 354175 156658 354184
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 150624 5228 150676 5234
rect 150624 5170 150676 5176
rect 150636 480 150664 5170
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 156512 9444 156564 9450
rect 156512 9386 156564 9392
rect 156524 3482 156552 9386
rect 156616 3670 156644 354175
rect 157340 352776 157392 352782
rect 157340 352718 157392 352724
rect 157352 16574 157380 352718
rect 160100 46232 160152 46238
rect 160100 46174 160152 46180
rect 157352 16546 157840 16574
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 156524 3454 156644 3482
rect 156616 480 156644 3454
rect 157812 480 157840 16546
rect 159364 10804 159416 10810
rect 159364 10746 159416 10752
rect 158904 7812 158956 7818
rect 158904 7754 158956 7760
rect 158916 480 158944 7754
rect 159376 3874 159404 10746
rect 159364 3868 159416 3874
rect 159364 3810 159416 3816
rect 160112 480 160140 46174
rect 162872 16574 162900 397054
rect 168380 394120 168432 394126
rect 168380 394062 168432 394068
rect 164240 392692 164292 392698
rect 164240 392634 164292 392640
rect 164252 16574 164280 392634
rect 162872 16546 163452 16574
rect 164252 16546 164464 16574
rect 162492 5296 162544 5302
rect 162492 5238 162544 5244
rect 161296 3664 161348 3670
rect 161296 3606 161348 3612
rect 161308 480 161336 3606
rect 162504 480 162532 5238
rect 163424 3482 163452 16546
rect 163504 15020 163556 15026
rect 163504 14962 163556 14968
rect 163516 3738 163544 14962
rect 163504 3732 163556 3738
rect 163504 3674 163556 3680
rect 163424 3454 163728 3482
rect 163700 480 163728 3454
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 167184 7880 167236 7886
rect 167184 7822 167236 7828
rect 166080 3868 166132 3874
rect 166080 3810 166132 3816
rect 166092 480 166120 3810
rect 167196 480 167224 7822
rect 168392 3398 168420 394062
rect 171152 16574 171180 398210
rect 184216 358766 184244 446150
rect 200764 445188 200816 445194
rect 200764 445130 200816 445136
rect 199384 445120 199436 445126
rect 199384 445062 199436 445068
rect 186964 444984 187016 444990
rect 186964 444926 187016 444932
rect 184940 391264 184992 391270
rect 184940 391206 184992 391212
rect 184204 358760 184256 358766
rect 184204 358702 184256 358708
rect 172518 352880 172574 352889
rect 172518 352815 172574 352824
rect 172532 16574 172560 352815
rect 182180 351348 182232 351354
rect 182180 351290 182232 351296
rect 180800 17264 180852 17270
rect 180800 17206 180852 17212
rect 180812 16574 180840 17206
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 180812 16546 181024 16574
rect 170770 7848 170826 7857
rect 170770 7783 170826 7792
rect 168472 3800 168524 3806
rect 168472 3742 168524 3748
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 168484 1986 168512 3742
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 168392 1958 168512 1986
rect 168392 480 168420 1958
rect 169588 480 169616 3334
rect 170784 480 170812 7783
rect 171980 480 172008 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 174266 9072 174322 9081
rect 174266 9007 174322 9016
rect 174280 480 174308 9007
rect 180248 6520 180300 6526
rect 180248 6462 180300 6468
rect 176660 6452 176712 6458
rect 176660 6394 176712 6400
rect 175462 3360 175518 3369
rect 175462 3295 175518 3304
rect 175476 480 175504 3295
rect 176672 480 176700 6394
rect 177856 4004 177908 4010
rect 177856 3946 177908 3952
rect 177868 480 177896 3946
rect 179052 3732 179104 3738
rect 179052 3674 179104 3680
rect 179064 480 179092 3674
rect 180260 480 180288 6462
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 351290
rect 183744 6588 183796 6594
rect 183744 6530 183796 6536
rect 183756 480 183784 6530
rect 184952 3398 184980 391206
rect 186976 267714 187004 444926
rect 191104 443284 191156 443290
rect 191104 443226 191156 443232
rect 188344 398404 188396 398410
rect 188344 398346 188396 398352
rect 187698 353016 187754 353025
rect 187698 352951 187754 352960
rect 186964 267708 187016 267714
rect 186964 267650 187016 267656
rect 187712 16574 187740 352951
rect 187712 16546 188292 16574
rect 187332 6656 187384 6662
rect 187332 6598 187384 6604
rect 185032 4072 185084 4078
rect 185032 4014 185084 4020
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 185044 2122 185072 4014
rect 186136 3392 186188 3398
rect 186136 3334 186188 3340
rect 184952 2094 185072 2122
rect 184952 480 184980 2094
rect 186148 480 186176 3334
rect 187344 480 187372 6598
rect 187700 5364 187752 5370
rect 187700 5306 187752 5312
rect 187712 3942 187740 5306
rect 187700 3936 187752 3942
rect 187700 3878 187752 3884
rect 188264 3482 188292 16546
rect 188356 6186 188384 398346
rect 189080 398336 189132 398342
rect 189080 398278 189132 398284
rect 189092 16574 189120 398278
rect 191116 241466 191144 443226
rect 198740 397180 198792 397186
rect 198740 397122 198792 397128
rect 191838 396944 191894 396953
rect 191838 396879 191894 396888
rect 191104 241460 191156 241466
rect 191104 241402 191156 241408
rect 191852 16574 191880 396879
rect 195980 394188 196032 394194
rect 195980 394130 196032 394136
rect 195992 16574 196020 394130
rect 189092 16546 189304 16574
rect 191852 16546 192064 16574
rect 195992 16546 196848 16574
rect 188344 6180 188396 6186
rect 188344 6122 188396 6128
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 190840 480 190868 3334
rect 192036 480 192064 16546
rect 195612 7948 195664 7954
rect 195612 7890 195664 7896
rect 194414 6216 194470 6225
rect 194414 6151 194470 6160
rect 193220 3936 193272 3942
rect 193220 3878 193272 3884
rect 193232 480 193260 3878
rect 194428 480 194456 6151
rect 195624 480 195652 7890
rect 196820 480 196848 16546
rect 197912 6180 197964 6186
rect 197912 6122 197964 6128
rect 197924 480 197952 6122
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 397122
rect 199396 164218 199424 445062
rect 199384 164212 199436 164218
rect 199384 164154 199436 164160
rect 200776 111790 200804 445130
rect 200868 411262 200896 446286
rect 202420 446276 202472 446282
rect 204350 446247 204406 446256
rect 202420 446218 202472 446224
rect 201958 446040 202014 446049
rect 201958 445975 202014 445984
rect 200856 411256 200908 411262
rect 200856 411198 200908 411204
rect 201972 352578 202000 445975
rect 202328 445256 202380 445262
rect 202328 445198 202380 445204
rect 202236 443896 202288 443902
rect 202236 443838 202288 443844
rect 202052 443624 202104 443630
rect 202052 443566 202104 443572
rect 201960 352572 202012 352578
rect 201960 352514 202012 352520
rect 202064 346390 202092 443566
rect 202142 442368 202198 442377
rect 202142 442303 202198 442312
rect 202052 346384 202104 346390
rect 202052 346326 202104 346332
rect 201500 177540 201552 177546
rect 201500 177482 201552 177488
rect 200764 111784 200816 111790
rect 200764 111726 200816 111732
rect 201408 5432 201460 5438
rect 201408 5374 201460 5380
rect 200304 4140 200356 4146
rect 200304 4082 200356 4088
rect 200316 480 200344 4082
rect 201420 3874 201448 5374
rect 201408 3868 201460 3874
rect 201408 3810 201460 3816
rect 201512 480 201540 177482
rect 202156 20670 202184 442303
rect 202248 59362 202276 443838
rect 202340 71738 202368 445198
rect 202432 85542 202460 446218
rect 204168 445800 204220 445806
rect 204168 445742 204220 445748
rect 203616 445324 203668 445330
rect 203616 445266 203668 445272
rect 203524 443828 203576 443834
rect 203524 443770 203576 443776
rect 202604 443760 202656 443766
rect 202604 443702 202656 443708
rect 203430 443728 203486 443737
rect 202510 442504 202566 442513
rect 202510 442439 202566 442448
rect 202524 97986 202552 442439
rect 202616 202842 202644 443702
rect 203430 443663 203486 443672
rect 202788 443556 202840 443562
rect 202788 443498 202840 443504
rect 202694 442640 202750 442649
rect 202694 442575 202750 442584
rect 202604 202836 202656 202842
rect 202604 202778 202656 202784
rect 202708 150414 202736 442575
rect 202800 293962 202828 443498
rect 202880 443352 202932 443358
rect 202880 443294 202932 443300
rect 202788 293956 202840 293962
rect 202788 293898 202840 293904
rect 202696 150408 202748 150414
rect 202696 150350 202748 150356
rect 202512 97980 202564 97986
rect 202512 97922 202564 97928
rect 202420 85536 202472 85542
rect 202420 85478 202472 85484
rect 202328 71732 202380 71738
rect 202328 71674 202380 71680
rect 202236 59356 202288 59362
rect 202236 59298 202288 59304
rect 202892 33114 202920 443294
rect 203444 443290 203472 443663
rect 203432 443284 203484 443290
rect 203432 443226 203484 443232
rect 202972 441516 203024 441522
rect 202972 441458 203024 441464
rect 202984 58682 203012 441458
rect 203064 177608 203116 177614
rect 203064 177550 203116 177556
rect 202972 58676 203024 58682
rect 202972 58618 203024 58624
rect 202880 33108 202932 33114
rect 202880 33050 202932 33056
rect 202144 20664 202196 20670
rect 202144 20606 202196 20612
rect 203076 16574 203104 177550
rect 203536 33046 203564 443770
rect 203628 215286 203656 445266
rect 204180 443698 204208 445742
rect 204364 443972 204392 446247
rect 204626 446176 204682 446185
rect 204626 446111 204682 446120
rect 204640 443972 204668 446111
rect 204916 445058 204944 446626
rect 209042 446584 209098 446593
rect 209042 446519 209098 446528
rect 206834 446448 206890 446457
rect 206834 446383 206890 446392
rect 206560 446140 206612 446146
rect 206560 446082 206612 446088
rect 204904 445052 204956 445058
rect 204904 444994 204956 445000
rect 205454 444816 205510 444825
rect 205454 444751 205510 444760
rect 205468 443972 205496 444751
rect 205730 444680 205786 444689
rect 205730 444615 205786 444624
rect 205744 443972 205772 444615
rect 206282 444544 206338 444553
rect 206282 444479 206338 444488
rect 206296 443972 206324 444479
rect 206572 443972 206600 446082
rect 206848 443972 206876 446383
rect 208216 446072 208268 446078
rect 208216 446014 208268 446020
rect 207110 444952 207166 444961
rect 207110 444887 207166 444896
rect 207124 443972 207152 444887
rect 207664 444644 207716 444650
rect 207664 444586 207716 444592
rect 207676 443972 207704 444586
rect 208228 443972 208256 446014
rect 208768 444372 208820 444378
rect 208768 444314 208820 444320
rect 208492 444100 208544 444106
rect 208492 444042 208544 444048
rect 208504 443972 208532 444042
rect 208780 443972 208808 444314
rect 209056 443972 209084 446519
rect 209320 444712 209372 444718
rect 209320 444654 209372 444660
rect 209332 443972 209360 444654
rect 209608 443972 209636 446655
rect 211252 446004 211304 446010
rect 211252 445946 211304 445952
rect 209872 445936 209924 445942
rect 209872 445878 209924 445884
rect 209884 443972 209912 445878
rect 210148 444848 210200 444854
rect 210148 444790 210200 444796
rect 210160 443972 210188 444790
rect 211264 443972 211292 445946
rect 211356 444786 211384 456758
rect 211528 455592 211580 455598
rect 211528 455534 211580 455540
rect 211436 455456 211488 455462
rect 211436 455398 211488 455404
rect 211448 446622 211476 455398
rect 211436 446616 211488 446622
rect 211436 446558 211488 446564
rect 211344 444780 211396 444786
rect 211344 444722 211396 444728
rect 211540 443972 211568 455534
rect 211816 449886 211844 487902
rect 215944 487688 215996 487694
rect 215944 487630 215996 487636
rect 214564 487620 214616 487626
rect 214564 487562 214616 487568
rect 213182 487520 213238 487529
rect 213182 487455 213238 487464
rect 213196 487422 213224 487455
rect 213184 487416 213236 487422
rect 213184 487358 213236 487364
rect 212448 487348 212500 487354
rect 212448 487290 212500 487296
rect 212460 486538 212488 487290
rect 212448 486532 212500 486538
rect 212448 486474 212500 486480
rect 212540 464364 212592 464370
rect 212540 464306 212592 464312
rect 211804 449880 211856 449886
rect 211804 449822 211856 449828
rect 212552 446758 212580 464306
rect 212724 463004 212776 463010
rect 212724 462946 212776 462952
rect 212632 446820 212684 446826
rect 212632 446762 212684 446768
rect 212356 446752 212408 446758
rect 212356 446694 212408 446700
rect 212540 446752 212592 446758
rect 212540 446694 212592 446700
rect 211804 446616 211856 446622
rect 211804 446558 211856 446564
rect 211816 443972 211844 446558
rect 212080 444780 212132 444786
rect 212080 444722 212132 444728
rect 212092 443972 212120 444722
rect 212368 443972 212396 446694
rect 212644 443972 212672 446762
rect 212736 443986 212764 462946
rect 212816 460216 212868 460222
rect 212816 460158 212868 460164
rect 212828 446622 212856 460158
rect 213196 459542 213224 487358
rect 214576 487257 214604 487562
rect 215956 487257 215984 487630
rect 214562 487248 214618 487257
rect 214562 487183 214618 487192
rect 215942 487248 215998 487257
rect 215942 487183 215998 487192
rect 214576 476066 214604 487183
rect 214564 476060 214616 476066
rect 214564 476002 214616 476008
rect 215956 471986 215984 487183
rect 218060 472660 218112 472666
rect 218060 472602 218112 472608
rect 215944 471980 215996 471986
rect 215944 471922 215996 471928
rect 217324 470620 217376 470626
rect 217324 470562 217376 470568
rect 216864 469940 216916 469946
rect 216864 469882 216916 469888
rect 216680 469872 216732 469878
rect 216680 469814 216732 469820
rect 213920 468580 213972 468586
rect 213920 468522 213972 468528
rect 213184 459536 213236 459542
rect 213184 459478 213236 459484
rect 213552 457496 213604 457502
rect 213552 457438 213604 457444
rect 213184 446752 213236 446758
rect 213184 446694 213236 446700
rect 212816 446616 212868 446622
rect 212816 446558 212868 446564
rect 213090 444136 213146 444145
rect 213090 444071 213146 444080
rect 212736 443958 212934 443986
rect 210332 443896 210384 443902
rect 207570 443864 207626 443873
rect 207414 443822 207570 443850
rect 210332 443838 210384 443844
rect 210884 443896 210936 443902
rect 211066 443864 211122 443873
rect 210884 443838 210936 443844
rect 207570 443799 207626 443808
rect 207966 443698 208164 443714
rect 204168 443692 204220 443698
rect 207966 443692 208176 443698
rect 207966 443686 208124 443692
rect 204168 443634 204220 443640
rect 208124 443634 208176 443640
rect 205086 443592 205142 443601
rect 204930 443550 205086 443578
rect 205086 443527 205142 443536
rect 205362 443456 205418 443465
rect 203904 443414 204102 443442
rect 205206 443414 205362 443442
rect 203904 443358 203932 443414
rect 206190 443456 206246 443465
rect 206034 443414 206190 443442
rect 205362 443391 205418 443400
rect 210344 443426 210372 443838
rect 210606 443456 210662 443465
rect 206190 443391 206246 443400
rect 210332 443420 210384 443426
rect 210450 443414 210606 443442
rect 210726 443426 210832 443442
rect 210896 443426 210924 443838
rect 211002 443822 211066 443850
rect 211066 443799 211122 443808
rect 211160 443828 211212 443834
rect 211160 443770 211212 443776
rect 211172 443494 211200 443770
rect 213104 443698 213132 444071
rect 213196 443972 213224 446694
rect 213460 446616 213512 446622
rect 213460 446558 213512 446564
rect 213472 443972 213500 446558
rect 213564 443986 213592 457438
rect 213932 446622 213960 468522
rect 215300 468512 215352 468518
rect 215300 468454 215352 468460
rect 214104 467152 214156 467158
rect 214104 467094 214156 467100
rect 214012 453552 214064 453558
rect 214012 453494 214064 453500
rect 213920 446616 213972 446622
rect 213920 446558 213972 446564
rect 213564 443958 213762 443986
rect 214024 443972 214052 453494
rect 214116 443986 214144 467094
rect 214196 464432 214248 464438
rect 214196 464374 214248 464380
rect 214208 444174 214236 464374
rect 214380 460284 214432 460290
rect 214380 460226 214432 460232
rect 214196 444168 214248 444174
rect 214196 444110 214248 444116
rect 214392 443986 214420 460226
rect 215116 446616 215168 446622
rect 215116 446558 215168 446564
rect 214840 444168 214892 444174
rect 214840 444110 214892 444116
rect 214116 443958 214314 443986
rect 214392 443958 214590 443986
rect 214852 443972 214880 444110
rect 215128 443972 215156 446558
rect 215312 444446 215340 468454
rect 215484 465724 215536 465730
rect 215484 465666 215536 465672
rect 215392 460352 215444 460358
rect 215392 460294 215444 460300
rect 215300 444440 215352 444446
rect 215300 444382 215352 444388
rect 215404 443972 215432 460294
rect 215496 444718 215524 465666
rect 215576 461712 215628 461718
rect 215576 461654 215628 461660
rect 215588 446622 215616 461654
rect 215668 454844 215720 454850
rect 215668 454786 215720 454792
rect 215576 446616 215628 446622
rect 215576 446558 215628 446564
rect 215484 444712 215536 444718
rect 215484 444654 215536 444660
rect 215680 443972 215708 454786
rect 216692 446622 216720 469814
rect 216772 461644 216824 461650
rect 216772 461586 216824 461592
rect 216220 446616 216272 446622
rect 216220 446558 216272 446564
rect 216680 446616 216732 446622
rect 216680 446558 216732 446564
rect 215944 444440 215996 444446
rect 215944 444382 215996 444388
rect 215956 443972 215984 444382
rect 216232 443972 216260 446558
rect 216496 444712 216548 444718
rect 216496 444654 216548 444660
rect 216588 444712 216640 444718
rect 216588 444654 216640 444660
rect 216508 443972 216536 444654
rect 216600 444106 216628 444654
rect 216588 444100 216640 444106
rect 216588 444042 216640 444048
rect 216680 444100 216732 444106
rect 216680 444042 216732 444048
rect 213092 443692 213144 443698
rect 213092 443634 213144 443640
rect 211160 443488 211212 443494
rect 211160 443430 211212 443436
rect 216692 443426 216720 444042
rect 216784 443972 216812 461586
rect 216876 444582 216904 469882
rect 216956 463072 217008 463078
rect 216956 463014 217008 463020
rect 216864 444576 216916 444582
rect 216864 444518 216916 444524
rect 216968 444514 216996 463014
rect 217048 461848 217100 461854
rect 217048 461790 217100 461796
rect 216956 444508 217008 444514
rect 216956 444450 217008 444456
rect 217060 443972 217088 461790
rect 217336 446826 217364 470562
rect 218072 447370 218100 472602
rect 218244 467288 218296 467294
rect 218244 467230 218296 467236
rect 218152 465792 218204 465798
rect 218152 465734 218204 465740
rect 218060 447364 218112 447370
rect 218060 447306 218112 447312
rect 217324 446820 217376 446826
rect 217324 446762 217376 446768
rect 217324 446616 217376 446622
rect 217324 446558 217376 446564
rect 217336 443972 217364 446558
rect 217600 444576 217652 444582
rect 217600 444518 217652 444524
rect 217414 444000 217470 444009
rect 217612 443972 217640 444518
rect 217876 444508 217928 444514
rect 217876 444450 217928 444456
rect 217888 443972 217916 444450
rect 218164 443972 218192 465734
rect 218256 447302 218284 467230
rect 218336 464500 218388 464506
rect 218336 464442 218388 464448
rect 218244 447296 218296 447302
rect 218244 447238 218296 447244
rect 218348 443986 218376 464442
rect 219532 453484 219584 453490
rect 219532 453426 219584 453432
rect 218704 450696 218756 450702
rect 218704 450638 218756 450644
rect 218348 443958 218454 443986
rect 218716 443972 218744 450638
rect 219072 447364 219124 447370
rect 219072 447306 219124 447312
rect 218796 447296 218848 447302
rect 218796 447238 218848 447244
rect 218808 443986 218836 447238
rect 219084 443986 219112 447306
rect 219440 444100 219492 444106
rect 219440 444042 219492 444048
rect 218808 443958 219006 443986
rect 219084 443958 219282 443986
rect 217414 443935 217470 443944
rect 217428 443737 217456 443935
rect 219346 443864 219402 443873
rect 219164 443828 219216 443834
rect 219346 443799 219402 443808
rect 219164 443770 219216 443776
rect 217414 443728 217470 443737
rect 217414 443663 217470 443672
rect 219176 443494 219204 443770
rect 219360 443630 219388 443799
rect 219348 443624 219400 443630
rect 219348 443566 219400 443572
rect 219164 443488 219216 443494
rect 219164 443430 219216 443436
rect 219452 443426 219480 444042
rect 219544 443972 219572 453426
rect 219636 443986 219664 487902
rect 219898 487792 219954 487801
rect 219898 487727 219954 487736
rect 219714 476776 219770 476785
rect 219714 476711 219770 476720
rect 219728 447134 219756 476711
rect 219912 460934 219940 487727
rect 220740 479534 220768 488407
rect 220728 479528 220780 479534
rect 220728 479470 220780 479476
rect 221096 475516 221148 475522
rect 221096 475458 221148 475464
rect 221108 460934 221136 475458
rect 224132 475448 224184 475454
rect 224132 475390 224184 475396
rect 224040 475380 224092 475386
rect 224040 475322 224092 475328
rect 221280 471300 221332 471306
rect 221280 471242 221332 471248
rect 221292 460934 221320 471242
rect 222660 463140 222712 463146
rect 222660 463082 222712 463088
rect 219912 460906 220216 460934
rect 221108 460906 221228 460934
rect 221292 460906 221596 460934
rect 219728 447106 219940 447134
rect 219912 443986 219940 447106
rect 220188 443986 220216 460906
rect 221004 452124 221056 452130
rect 221004 452066 221056 452072
rect 221016 447302 221044 452066
rect 221096 450764 221148 450770
rect 221096 450706 221148 450712
rect 221004 447296 221056 447302
rect 221004 447238 221056 447244
rect 220636 446480 220688 446486
rect 220636 446422 220688 446428
rect 220450 444000 220506 444009
rect 219636 443958 219834 443986
rect 219912 443958 220110 443986
rect 220188 443958 220386 443986
rect 220648 443972 220676 446422
rect 220912 446412 220964 446418
rect 220912 446354 220964 446360
rect 220924 443972 220952 446354
rect 221108 443986 221136 450706
rect 221200 447134 221228 460906
rect 221200 447106 221320 447134
rect 221292 443986 221320 447106
rect 221568 443986 221596 460906
rect 222292 453416 222344 453422
rect 222292 453358 222344 453364
rect 221832 447296 221884 447302
rect 221832 447238 221884 447244
rect 221844 443986 221872 447238
rect 221108 443958 221214 443986
rect 221292 443958 221490 443986
rect 221568 443958 221766 443986
rect 221844 443958 222042 443986
rect 222304 443972 222332 453358
rect 222384 452056 222436 452062
rect 222384 451998 222436 452004
rect 222396 445058 222424 451998
rect 222568 447908 222620 447914
rect 222568 447850 222620 447856
rect 222580 446418 222608 447850
rect 222568 446412 222620 446418
rect 222568 446354 222620 446360
rect 222384 445052 222436 445058
rect 222384 444994 222436 445000
rect 222476 444032 222528 444038
rect 222476 443974 222528 443980
rect 220450 443935 220506 443944
rect 220464 443494 220492 443935
rect 222488 443562 222516 443974
rect 222580 443972 222608 446354
rect 222672 443986 222700 463082
rect 224052 460934 224080 475322
rect 223684 460906 224080 460934
rect 224144 460934 224172 475390
rect 225604 461780 225656 461786
rect 225604 461722 225656 461728
rect 224144 460906 224356 460934
rect 223212 456272 223264 456278
rect 223212 456214 223264 456220
rect 223224 448526 223252 456214
rect 223580 453348 223632 453354
rect 223580 453290 223632 453296
rect 223212 448520 223264 448526
rect 223212 448462 223264 448468
rect 222936 445052 222988 445058
rect 222936 444994 222988 445000
rect 222948 443986 222976 444994
rect 223224 443986 223252 448462
rect 223592 444258 223620 453290
rect 223684 444378 223712 460906
rect 224040 455524 224092 455530
rect 224040 455466 224092 455472
rect 224052 455394 224080 455466
rect 223764 455388 223816 455394
rect 223764 455330 223816 455336
rect 224040 455388 224092 455394
rect 224040 455330 224092 455336
rect 223776 447134 223804 455330
rect 223776 447106 224080 447134
rect 223672 444372 223724 444378
rect 223672 444314 223724 444320
rect 223592 444230 223804 444258
rect 223672 444100 223724 444106
rect 223672 444042 223724 444048
rect 222672 443958 222870 443986
rect 222948 443958 223146 443986
rect 223224 443958 223422 443986
rect 223684 443972 223712 444042
rect 223776 443986 223804 444230
rect 224052 443986 224080 447106
rect 224328 443986 224356 460906
rect 224960 457564 225012 457570
rect 224960 457506 225012 457512
rect 224972 455734 225000 457506
rect 224960 455728 225012 455734
rect 224960 455670 225012 455676
rect 225420 455728 225472 455734
rect 225420 455670 225472 455676
rect 225144 451920 225196 451926
rect 225144 451862 225196 451868
rect 224776 450628 224828 450634
rect 224776 450570 224828 450576
rect 223776 443958 223974 443986
rect 224052 443958 224250 443986
rect 224328 443958 224526 443986
rect 224788 443972 224816 450570
rect 225156 447302 225184 451862
rect 225328 450560 225380 450566
rect 225328 450502 225380 450508
rect 225144 447296 225196 447302
rect 225144 447238 225196 447244
rect 225052 446820 225104 446826
rect 225052 446762 225104 446768
rect 225064 443972 225092 446762
rect 225340 443972 225368 450502
rect 225432 447370 225460 455670
rect 225512 454708 225564 454714
rect 225512 454650 225564 454656
rect 225420 447364 225472 447370
rect 225420 447306 225472 447312
rect 225524 443986 225552 454650
rect 225616 446826 225644 461722
rect 226260 451926 226288 488407
rect 226984 462392 227036 462398
rect 226984 462334 227036 462340
rect 226616 454776 226668 454782
rect 226616 454718 226668 454724
rect 226248 451920 226300 451926
rect 226248 451862 226300 451868
rect 225696 447364 225748 447370
rect 225696 447306 225748 447312
rect 225604 446820 225656 446826
rect 225604 446762 225656 446768
rect 225708 443986 225736 447306
rect 225972 447296 226024 447302
rect 225972 447238 226024 447244
rect 225984 443986 226012 447238
rect 226628 443986 226656 454718
rect 226892 451988 226944 451994
rect 226892 451930 226944 451936
rect 226708 446888 226760 446894
rect 226708 446830 226760 446836
rect 225524 443958 225630 443986
rect 225708 443958 225906 443986
rect 225984 443958 226182 443986
rect 226458 443958 226656 443986
rect 226720 443972 226748 446830
rect 226904 443986 226932 451930
rect 226996 444514 227024 462334
rect 227076 457632 227128 457638
rect 227076 457574 227128 457580
rect 227088 446894 227116 457574
rect 231124 456884 231176 456890
rect 231124 456826 231176 456832
rect 228546 454064 228602 454073
rect 228546 453999 228602 454008
rect 227260 447840 227312 447846
rect 227260 447782 227312 447788
rect 227076 446888 227128 446894
rect 227076 446830 227128 446836
rect 226984 444508 227036 444514
rect 226984 444450 227036 444456
rect 226904 443958 227010 443986
rect 227272 443972 227300 447782
rect 228364 446344 228416 446350
rect 228364 446286 228416 446292
rect 227812 444916 227864 444922
rect 227812 444858 227864 444864
rect 227536 444508 227588 444514
rect 227536 444450 227588 444456
rect 227548 443972 227576 444450
rect 227824 443972 227852 444858
rect 228376 443986 228404 446286
rect 228560 445398 228588 453999
rect 229468 446752 229520 446758
rect 229468 446694 229520 446700
rect 229008 446616 229060 446622
rect 229008 446558 229060 446564
rect 229020 446457 229048 446558
rect 229100 446480 229152 446486
rect 229006 446448 229062 446457
rect 229100 446422 229152 446428
rect 229006 446383 229062 446392
rect 229112 446321 229140 446422
rect 229098 446312 229154 446321
rect 229098 446247 229154 446256
rect 229192 446208 229244 446214
rect 229192 446150 229244 446156
rect 228548 445392 228600 445398
rect 228548 445334 228600 445340
rect 228560 443986 228588 445334
rect 228376 443972 228496 443986
rect 228390 443958 228496 443972
rect 228560 443958 228666 443986
rect 229204 443972 229232 446150
rect 229480 445466 229508 446694
rect 230848 446548 230900 446554
rect 230848 446490 230900 446496
rect 229652 446412 229704 446418
rect 229652 446354 229704 446360
rect 229744 446412 229796 446418
rect 229744 446354 229796 446360
rect 229468 445460 229520 445466
rect 229468 445402 229520 445408
rect 229480 443972 229508 445402
rect 229664 445058 229692 446354
rect 229756 446185 229784 446354
rect 229742 446176 229798 446185
rect 229742 446111 229798 446120
rect 230020 445868 230072 445874
rect 230020 445810 230072 445816
rect 229652 445052 229704 445058
rect 229652 444994 229704 445000
rect 230032 443972 230060 445810
rect 230296 444984 230348 444990
rect 230296 444926 230348 444932
rect 230308 444446 230336 444926
rect 230296 444440 230348 444446
rect 230296 444382 230348 444388
rect 230308 443972 230336 444382
rect 230860 443972 230888 446490
rect 231136 445330 231164 456826
rect 231780 447846 231808 488446
rect 235630 487928 235686 487937
rect 235630 487863 235686 487872
rect 235644 487830 235672 487863
rect 235632 487824 235684 487830
rect 235632 487766 235684 487772
rect 235908 487824 235960 487830
rect 235908 487766 235960 487772
rect 232136 457224 232188 457230
rect 232136 457166 232188 457172
rect 231768 447840 231820 447846
rect 231768 447782 231820 447788
rect 232148 447134 232176 457166
rect 232596 457020 232648 457026
rect 232596 456962 232648 456968
rect 231964 447106 232176 447134
rect 231400 446684 231452 446690
rect 231400 446626 231452 446632
rect 231124 445324 231176 445330
rect 231124 445266 231176 445272
rect 231136 443972 231164 445266
rect 231412 443972 231440 446626
rect 231964 445126 231992 447106
rect 232228 445800 232280 445806
rect 232228 445742 232280 445748
rect 231952 445120 232004 445126
rect 231952 445062 232004 445068
rect 231504 443970 231702 443986
rect 231964 443972 231992 445062
rect 232240 443972 232268 445742
rect 232608 445194 232636 456962
rect 235920 447914 235948 487766
rect 240140 481024 240192 481030
rect 240140 480966 240192 480972
rect 236000 480956 236052 480962
rect 236000 480898 236052 480904
rect 235908 447908 235960 447914
rect 235908 447850 235960 447856
rect 236012 447370 236040 480898
rect 239956 479596 240008 479602
rect 239956 479538 240008 479544
rect 236368 476808 236420 476814
rect 236368 476750 236420 476756
rect 236184 467220 236236 467226
rect 236184 467162 236236 467168
rect 236000 447364 236052 447370
rect 236000 447306 236052 447312
rect 235538 446856 235594 446865
rect 235538 446791 235594 446800
rect 233606 446312 233662 446321
rect 233056 446276 233108 446282
rect 233606 446247 233662 446256
rect 233056 446218 233108 446224
rect 232596 445188 232648 445194
rect 232596 445130 232648 445136
rect 232780 445188 232832 445194
rect 232780 445130 232832 445136
rect 232792 443972 232820 445130
rect 233068 443972 233096 446218
rect 233620 445262 233648 446247
rect 234710 446040 234766 446049
rect 234710 445975 234766 445984
rect 233608 445256 233660 445262
rect 233608 445198 233660 445204
rect 233620 443972 233648 445198
rect 234436 444916 234488 444922
rect 234436 444858 234488 444864
rect 231492 443964 231702 443970
rect 228468 443834 228496 443958
rect 231544 443958 231702 443964
rect 231492 443906 231544 443912
rect 228732 443896 228784 443902
rect 232318 443864 232374 443873
rect 228784 443844 228942 443850
rect 228732 443838 228942 443844
rect 222752 443828 222804 443834
rect 222752 443770 222804 443776
rect 228456 443828 228508 443834
rect 228744 443822 228942 443838
rect 233238 443864 233294 443873
rect 232374 443822 232530 443850
rect 232318 443799 232374 443808
rect 233294 443822 233358 443850
rect 233238 443799 233294 443808
rect 228456 443770 228508 443776
rect 222764 443698 222792 443770
rect 229560 443760 229612 443766
rect 234448 443714 234476 444858
rect 234724 443972 234752 445975
rect 235262 445088 235318 445097
rect 235262 445023 235318 445032
rect 235276 443972 235304 445023
rect 235552 443972 235580 446791
rect 236196 443986 236224 467162
rect 236276 463140 236328 463146
rect 236276 463082 236328 463088
rect 236288 447302 236316 463082
rect 236276 447296 236328 447302
rect 236276 447238 236328 447244
rect 236118 443958 236224 443986
rect 236380 443972 236408 476750
rect 238116 475448 238168 475454
rect 238116 475390 238168 475396
rect 238024 474020 238076 474026
rect 238024 473962 238076 473968
rect 237932 458924 237984 458930
rect 237932 458866 237984 458872
rect 237840 458312 237892 458318
rect 237840 458254 237892 458260
rect 237564 455796 237616 455802
rect 237564 455738 237616 455744
rect 237472 448452 237524 448458
rect 237472 448394 237524 448400
rect 236460 447364 236512 447370
rect 236460 447306 236512 447312
rect 236472 443986 236500 447306
rect 236736 447296 236788 447302
rect 236736 447238 236788 447244
rect 236748 443986 236776 447238
rect 237196 444984 237248 444990
rect 237196 444926 237248 444932
rect 236472 443958 236670 443986
rect 236748 443958 236946 443986
rect 237208 443972 237236 444926
rect 237484 443972 237512 448394
rect 237576 445330 237604 455738
rect 237746 446176 237802 446185
rect 237746 446111 237802 446120
rect 237564 445324 237616 445330
rect 237564 445266 237616 445272
rect 237760 443972 237788 446111
rect 237852 443986 237880 458254
rect 237944 446554 237972 458866
rect 238036 448458 238064 473962
rect 238128 459406 238156 475390
rect 239968 474706 239996 479538
rect 240048 478236 240100 478242
rect 240048 478178 240100 478184
rect 238760 474700 238812 474706
rect 238760 474642 238812 474648
rect 239956 474700 240008 474706
rect 239956 474642 240008 474648
rect 238208 471300 238260 471306
rect 238208 471242 238260 471248
rect 238220 459474 238248 471242
rect 238208 459468 238260 459474
rect 238208 459410 238260 459416
rect 238116 459400 238168 459406
rect 238116 459342 238168 459348
rect 238128 458318 238156 459342
rect 238220 458930 238248 459410
rect 238208 458924 238260 458930
rect 238208 458866 238260 458872
rect 238116 458312 238168 458318
rect 238116 458254 238168 458260
rect 238024 448452 238076 448458
rect 238024 448394 238076 448400
rect 237932 446548 237984 446554
rect 237932 446490 237984 446496
rect 238576 446548 238628 446554
rect 238576 446490 238628 446496
rect 238300 445324 238352 445330
rect 238300 445266 238352 445272
rect 237852 443958 238050 443986
rect 238312 443972 238340 445266
rect 238588 443972 238616 446490
rect 238772 445466 238800 474642
rect 240060 473346 240088 478178
rect 240152 477494 240180 480966
rect 240140 477488 240192 477494
rect 240140 477430 240192 477436
rect 239128 473340 239180 473346
rect 239128 473282 239180 473288
rect 240048 473340 240100 473346
rect 240048 473282 240100 473288
rect 239036 455932 239088 455938
rect 239036 455874 239088 455880
rect 238944 455864 238996 455870
rect 238944 455806 238996 455812
rect 238956 446554 238984 455806
rect 238944 446548 238996 446554
rect 238944 446490 238996 446496
rect 238760 445460 238812 445466
rect 238760 445402 238812 445408
rect 239048 443986 239076 455874
rect 238878 443958 239076 443986
rect 239140 443972 239168 473282
rect 239956 446548 240008 446554
rect 239956 446490 240008 446496
rect 239680 445460 239732 445466
rect 239680 445402 239732 445408
rect 239404 445120 239456 445126
rect 239404 445062 239456 445068
rect 239416 443972 239444 445062
rect 239692 443972 239720 445402
rect 239968 443972 239996 446490
rect 240152 443986 240180 477430
rect 240796 452606 240824 489126
rect 242900 488776 242952 488782
rect 242900 488718 242952 488724
rect 241426 487928 241482 487937
rect 241426 487863 241482 487872
rect 241440 487830 241468 487863
rect 241428 487824 241480 487830
rect 241428 487766 241480 487772
rect 241440 487218 241468 487766
rect 241428 487212 241480 487218
rect 241428 487154 241480 487160
rect 240876 478168 240928 478174
rect 240876 478110 240928 478116
rect 240784 452600 240836 452606
rect 240784 452542 240836 452548
rect 240324 451308 240376 451314
rect 240324 451250 240376 451256
rect 240336 444310 240364 451250
rect 240692 449948 240744 449954
rect 240692 449890 240744 449896
rect 240324 444304 240376 444310
rect 240324 444246 240376 444252
rect 240704 443986 240732 449890
rect 240796 444394 240824 452542
rect 240888 451246 240916 478110
rect 241440 472734 241468 487154
rect 241520 486464 241572 486470
rect 241520 486406 241572 486412
rect 241532 484362 241560 486406
rect 241520 484356 241572 484362
rect 241520 484298 241572 484304
rect 241428 472728 241480 472734
rect 241428 472670 241480 472676
rect 240876 451240 240928 451246
rect 240876 451182 240928 451188
rect 240888 449954 240916 451182
rect 240876 449948 240928 449954
rect 240876 449890 240928 449896
rect 241532 446554 241560 484298
rect 242808 482384 242860 482390
rect 242808 482326 242860 482332
rect 241888 478848 241940 478854
rect 241888 478790 241940 478796
rect 241900 478038 241928 478790
rect 242820 478038 242848 482326
rect 241888 478032 241940 478038
rect 241888 477974 241940 477980
rect 242808 478032 242860 478038
rect 242808 477974 242860 477980
rect 241796 457292 241848 457298
rect 241796 457234 241848 457240
rect 241704 456952 241756 456958
rect 241704 456894 241756 456900
rect 241716 451110 241744 456894
rect 241704 451104 241756 451110
rect 241704 451046 241756 451052
rect 241520 446548 241572 446554
rect 241520 446490 241572 446496
rect 241612 446276 241664 446282
rect 241612 446218 241664 446224
rect 240796 444366 241192 444394
rect 241060 444304 241112 444310
rect 241060 444246 241112 444252
rect 240152 443958 240258 443986
rect 240704 443958 240810 443986
rect 241072 443972 241100 444246
rect 241164 443986 241192 444366
rect 241164 443958 241362 443986
rect 241624 443972 241652 446218
rect 241808 445262 241836 457234
rect 241796 445256 241848 445262
rect 241796 445198 241848 445204
rect 241900 443972 241928 477974
rect 241980 451104 242032 451110
rect 241980 451046 242032 451052
rect 241992 443986 242020 451046
rect 242440 446548 242492 446554
rect 242440 446490 242492 446496
rect 241992 443958 242190 443986
rect 242452 443972 242480 446490
rect 242912 446350 242940 488718
rect 244556 487892 244608 487898
rect 244556 487834 244608 487840
rect 244568 487354 244596 487834
rect 250442 487520 250498 487529
rect 250442 487455 250498 487464
rect 250456 487422 250484 487455
rect 250444 487416 250496 487422
rect 245566 487384 245622 487393
rect 244556 487348 244608 487354
rect 250444 487358 250496 487364
rect 251088 487416 251140 487422
rect 251088 487358 251140 487364
rect 245566 487319 245568 487328
rect 244556 487290 244608 487296
rect 245620 487319 245622 487328
rect 245568 487290 245620 487296
rect 244924 486464 244976 486470
rect 244924 486406 244976 486412
rect 243544 481092 243596 481098
rect 243544 481034 243596 481040
rect 243556 473346 243584 481034
rect 244280 479528 244332 479534
rect 244280 479470 244332 479476
rect 243084 473340 243136 473346
rect 243084 473282 243136 473288
rect 243544 473340 243596 473346
rect 243544 473282 243596 473288
rect 242992 457088 243044 457094
rect 242992 457030 243044 457036
rect 242900 446344 242952 446350
rect 242900 446286 242952 446292
rect 242716 445256 242768 445262
rect 242716 445198 242768 445204
rect 242728 443972 242756 445198
rect 243004 443972 243032 457030
rect 243096 445466 243124 473282
rect 244292 460934 244320 479470
rect 244936 460934 244964 486406
rect 245580 477494 245608 487290
rect 247684 486532 247736 486538
rect 247684 486474 247736 486480
rect 246120 482316 246172 482322
rect 246120 482258 246172 482264
rect 246132 480254 246160 482258
rect 245856 480226 246160 480254
rect 245856 478854 245884 480226
rect 245844 478848 245896 478854
rect 245844 478790 245896 478796
rect 245568 477488 245620 477494
rect 245568 477430 245620 477436
rect 245856 460934 245884 478790
rect 247696 474706 247724 486474
rect 250352 482316 250404 482322
rect 250352 482258 250404 482264
rect 249800 477488 249852 477494
rect 249800 477430 249852 477436
rect 249156 476808 249208 476814
rect 249156 476750 249208 476756
rect 249064 475380 249116 475386
rect 249064 475322 249116 475328
rect 247040 474700 247092 474706
rect 247040 474642 247092 474648
rect 247684 474700 247736 474706
rect 247684 474642 247736 474648
rect 247052 460934 247080 474642
rect 248696 472728 248748 472734
rect 248696 472670 248748 472676
rect 244292 460906 244412 460934
rect 244936 460906 245056 460934
rect 245856 460906 246160 460934
rect 247052 460906 247172 460934
rect 243636 457156 243688 457162
rect 243636 457098 243688 457104
rect 243544 446344 243596 446350
rect 243544 446286 243596 446292
rect 243084 445460 243136 445466
rect 243084 445402 243136 445408
rect 243556 443972 243584 446286
rect 243648 443986 243676 457098
rect 244384 449894 244412 460906
rect 244740 456000 244792 456006
rect 244740 455942 244792 455948
rect 244384 449866 244504 449894
rect 244372 446548 244424 446554
rect 244372 446490 244424 446496
rect 244096 445460 244148 445466
rect 244096 445402 244148 445408
rect 243648 443958 243846 443986
rect 244108 443972 244136 445402
rect 244384 443972 244412 446490
rect 244476 443986 244504 449866
rect 244752 443986 244780 455942
rect 245028 449818 245056 460906
rect 245752 451920 245804 451926
rect 245752 451862 245804 451868
rect 245016 449812 245068 449818
rect 245016 449754 245068 449760
rect 245028 443986 245056 449754
rect 245474 445632 245530 445641
rect 245474 445567 245530 445576
rect 244476 443958 244674 443986
rect 244752 443958 244950 443986
rect 245028 443958 245226 443986
rect 245488 443972 245516 445567
rect 245764 443972 245792 451862
rect 246132 443986 246160 460906
rect 246304 458924 246356 458930
rect 246304 458866 246356 458872
rect 246316 446554 246344 458866
rect 247144 449894 247172 460906
rect 248604 453348 248656 453354
rect 248604 453290 248656 453296
rect 248052 451920 248104 451926
rect 248052 451862 248104 451868
rect 247144 449866 247264 449894
rect 246856 447840 246908 447846
rect 246856 447782 246908 447788
rect 246304 446548 246356 446554
rect 246304 446490 246356 446496
rect 246132 443958 246330 443986
rect 246868 443972 246896 447782
rect 247132 446684 247184 446690
rect 247132 446626 247184 446632
rect 247144 443972 247172 446626
rect 247236 443986 247264 449866
rect 247960 447908 248012 447914
rect 247960 447850 248012 447856
rect 247684 447160 247736 447166
rect 247684 447102 247736 447108
rect 247500 446140 247552 446146
rect 247500 446082 247552 446088
rect 247512 444145 247540 446082
rect 247498 444136 247554 444145
rect 247498 444071 247554 444080
rect 247236 443958 247434 443986
rect 247696 443972 247724 447102
rect 247972 443972 248000 447850
rect 248064 443986 248092 451862
rect 248512 449880 248564 449886
rect 248512 449822 248564 449828
rect 248524 449478 248552 449822
rect 248512 449472 248564 449478
rect 248512 449414 248564 449420
rect 248064 443958 248262 443986
rect 248524 443972 248552 449414
rect 248616 443986 248644 453290
rect 248708 449894 248736 472670
rect 248972 459536 249024 459542
rect 248972 459478 249024 459484
rect 248708 449866 248920 449894
rect 248892 443986 248920 449866
rect 248984 445398 249012 459478
rect 249076 449478 249104 475322
rect 249168 459542 249196 476750
rect 249812 460934 249840 477430
rect 250364 476066 250392 482258
rect 251100 476218 251128 487358
rect 261484 485104 261536 485110
rect 261484 485046 261536 485052
rect 261576 485104 261628 485110
rect 261576 485046 261628 485052
rect 251640 479528 251692 479534
rect 251640 479470 251692 479476
rect 251100 476190 251220 476218
rect 250352 476060 250404 476066
rect 250352 476002 250404 476008
rect 250364 460934 250392 476002
rect 249812 460906 249932 460934
rect 250364 460906 250576 460934
rect 249156 459536 249208 459542
rect 249156 459478 249208 459484
rect 249904 449894 249932 460906
rect 250076 456068 250128 456074
rect 250076 456010 250128 456016
rect 249904 449866 250024 449894
rect 249064 449472 249116 449478
rect 249064 449414 249116 449420
rect 249892 445800 249944 445806
rect 249892 445742 249944 445748
rect 248972 445392 249024 445398
rect 248972 445334 249024 445340
rect 249616 445392 249668 445398
rect 249616 445334 249668 445340
rect 248616 443958 248814 443986
rect 248892 443958 249090 443986
rect 249628 443972 249656 445334
rect 249904 443972 249932 445742
rect 249996 443986 250024 449866
rect 250088 445602 250116 456010
rect 250442 445768 250498 445777
rect 250442 445703 250498 445712
rect 250076 445596 250128 445602
rect 250076 445538 250128 445544
rect 249996 443958 250194 443986
rect 250456 443972 250484 445703
rect 250548 443986 250576 460906
rect 250996 445596 251048 445602
rect 250996 445538 251048 445544
rect 250548 443958 250746 443986
rect 251008 443972 251036 445538
rect 251192 443986 251220 476190
rect 251652 471986 251680 479470
rect 251640 471980 251692 471986
rect 251640 471922 251692 471928
rect 251546 444408 251602 444417
rect 251546 444343 251602 444352
rect 251192 443958 251298 443986
rect 251560 443972 251588 444343
rect 251652 443986 251680 471922
rect 261208 469192 261260 469198
rect 261208 469134 261260 469140
rect 261220 468926 261248 469134
rect 261208 468920 261260 468926
rect 261208 468862 261260 468868
rect 260932 458856 260984 458862
rect 260932 458798 260984 458804
rect 260196 458516 260248 458522
rect 260196 458458 260248 458464
rect 254584 458312 254636 458318
rect 254584 458254 254636 458260
rect 254492 454776 254544 454782
rect 254492 454718 254544 454724
rect 252560 454708 252612 454714
rect 252560 454650 252612 454656
rect 252376 449336 252428 449342
rect 252376 449278 252428 449284
rect 252100 447840 252152 447846
rect 252100 447782 252152 447788
rect 251732 446616 251784 446622
rect 251732 446558 251784 446564
rect 251744 446049 251772 446558
rect 251824 446072 251876 446078
rect 251730 446040 251786 446049
rect 251824 446014 251876 446020
rect 251730 445975 251786 445984
rect 251836 445913 251864 446014
rect 251822 445904 251878 445913
rect 251822 445839 251878 445848
rect 251652 443958 251850 443986
rect 252112 443972 252140 447782
rect 252388 443972 252416 449278
rect 252572 443986 252600 454650
rect 253480 449472 253532 449478
rect 253480 449414 253532 449420
rect 252926 449168 252982 449177
rect 252926 449103 252982 449112
rect 252572 443958 252678 443986
rect 252940 443972 252968 449103
rect 253204 445868 253256 445874
rect 253204 445810 253256 445816
rect 253216 443972 253244 445810
rect 253492 443972 253520 449414
rect 254030 449304 254086 449313
rect 254030 449239 254086 449248
rect 254308 449268 254360 449274
rect 253756 449200 253808 449206
rect 253756 449142 253808 449148
rect 253768 443972 253796 449142
rect 254044 443972 254072 449239
rect 254308 449210 254360 449216
rect 254320 443972 254348 449210
rect 254400 446548 254452 446554
rect 254400 446490 254452 446496
rect 254412 443986 254440 446490
rect 254504 444122 254532 454718
rect 254596 445806 254624 458254
rect 258080 456204 258132 456210
rect 258080 456146 258132 456152
rect 255780 456136 255832 456142
rect 255780 456078 255832 456084
rect 255688 449676 255740 449682
rect 255688 449618 255740 449624
rect 255136 449540 255188 449546
rect 255136 449482 255188 449488
rect 254584 445800 254636 445806
rect 254584 445742 254636 445748
rect 254504 444094 254716 444122
rect 254688 443986 254716 444094
rect 254412 443958 254610 443986
rect 254688 443958 254886 443986
rect 255148 443972 255176 449482
rect 255412 446072 255464 446078
rect 255412 446014 255464 446020
rect 255424 443972 255452 446014
rect 255700 443972 255728 449618
rect 255792 443986 255820 456078
rect 257896 449812 257948 449818
rect 257896 449754 257948 449760
rect 257344 449608 257396 449614
rect 257344 449550 257396 449556
rect 256240 449404 256292 449410
rect 256240 449346 256292 449352
rect 255792 443958 255990 443986
rect 256252 443972 256280 449346
rect 256792 446616 256844 446622
rect 256792 446558 256844 446564
rect 256804 443972 256832 446558
rect 257356 443972 257384 449550
rect 257436 446276 257488 446282
rect 257436 446218 257488 446224
rect 249156 443896 249208 443902
rect 234894 443864 234950 443873
rect 234950 443822 235014 443850
rect 249156 443838 249208 443844
rect 250812 443896 250864 443902
rect 250812 443838 250864 443844
rect 243176 443828 243228 443834
rect 234894 443799 234950 443808
rect 243176 443770 243228 443776
rect 235908 443760 235960 443766
rect 229612 443708 229770 443714
rect 229560 443702 229770 443708
rect 222752 443692 222804 443698
rect 229572 443686 229770 443702
rect 234264 443700 234476 443714
rect 235842 443708 235908 443714
rect 235842 443702 235960 443708
rect 234264 443698 234462 443700
rect 234252 443692 234462 443698
rect 222752 443634 222804 443640
rect 234304 443686 234462 443692
rect 235842 443686 235948 443702
rect 234252 443634 234304 443640
rect 230480 443624 230532 443630
rect 230532 443572 230598 443578
rect 230480 443566 230598 443572
rect 222476 443556 222528 443562
rect 230492 443550 230598 443566
rect 233988 443562 234186 443578
rect 233976 443556 234186 443562
rect 222476 443498 222528 443504
rect 234028 443550 234186 443556
rect 240416 443556 240468 443562
rect 233976 443498 234028 443504
rect 240416 443498 240468 443504
rect 220452 443488 220504 443494
rect 220452 443430 220504 443436
rect 227916 443426 228114 443442
rect 233712 443426 233910 443442
rect 240428 443426 240456 443498
rect 240534 443426 240732 443442
rect 243188 443426 243216 443770
rect 246606 443698 246804 443714
rect 246606 443692 246816 443698
rect 246606 443686 246764 443692
rect 246764 443634 246816 443640
rect 248880 443624 248932 443630
rect 248880 443566 248932 443572
rect 243452 443488 243504 443494
rect 243294 443436 243452 443442
rect 246212 443488 246264 443494
rect 243294 443430 243504 443436
rect 246054 443436 246212 443442
rect 246054 443430 246264 443436
rect 210726 443420 210844 443426
rect 210726 443414 210792 443420
rect 210606 443391 210662 443400
rect 210332 443362 210384 443368
rect 210792 443362 210844 443368
rect 210884 443420 210936 443426
rect 210884 443362 210936 443368
rect 216680 443420 216732 443426
rect 216680 443362 216732 443368
rect 219440 443420 219492 443426
rect 219440 443362 219492 443368
rect 227904 443420 228114 443426
rect 227956 443414 228114 443420
rect 233700 443420 233910 443426
rect 227904 443362 227956 443368
rect 233752 443414 233910 443420
rect 240416 443420 240468 443426
rect 233700 443362 233752 443368
rect 240534 443420 240744 443426
rect 240534 443414 240692 443420
rect 240416 443362 240468 443368
rect 240692 443362 240744 443368
rect 243176 443420 243228 443426
rect 243294 443414 243492 443430
rect 246054 443414 246252 443430
rect 248892 443426 248920 443566
rect 248972 443556 249024 443562
rect 248972 443498 249024 443504
rect 248984 443426 249012 443498
rect 249168 443426 249196 443838
rect 249366 443426 249564 443442
rect 250824 443426 250852 443838
rect 250904 443828 250956 443834
rect 250904 443770 250956 443776
rect 251088 443828 251140 443834
rect 251088 443770 251140 443776
rect 251732 443828 251784 443834
rect 251732 443770 251784 443776
rect 250916 443426 250944 443770
rect 251100 443698 251128 443770
rect 251088 443692 251140 443698
rect 251088 443634 251140 443640
rect 251180 443692 251232 443698
rect 251180 443634 251232 443640
rect 251192 443494 251220 443634
rect 251180 443488 251232 443494
rect 251180 443430 251232 443436
rect 251744 443426 251772 443770
rect 257448 443698 257476 446218
rect 257620 446140 257672 446146
rect 257620 446082 257672 446088
rect 257632 443972 257660 446082
rect 257908 443972 257936 449754
rect 258092 443986 258120 456146
rect 259828 450560 259880 450566
rect 259828 450502 259880 450508
rect 259552 449880 259604 449886
rect 259552 449822 259604 449828
rect 258632 449744 258684 449750
rect 258632 449686 258684 449692
rect 258448 446412 258500 446418
rect 258448 446354 258500 446360
rect 258460 445641 258488 446354
rect 258446 445632 258502 445641
rect 258446 445567 258502 445576
rect 258644 443986 258672 449686
rect 259000 449064 259052 449070
rect 259000 449006 259052 449012
rect 258092 443958 258198 443986
rect 258474 443958 258672 443986
rect 259012 443972 259040 449006
rect 259564 443972 259592 449822
rect 259840 443972 259868 450502
rect 260104 448996 260156 449002
rect 260104 448938 260156 448944
rect 260116 443972 260144 448938
rect 260208 443986 260236 458458
rect 260656 449132 260708 449138
rect 260656 449074 260708 449080
rect 260208 443958 260406 443986
rect 260668 443972 260696 449074
rect 260840 446480 260892 446486
rect 260840 446422 260892 446428
rect 260852 446185 260880 446422
rect 260838 446176 260894 446185
rect 260838 446111 260894 446120
rect 260944 443972 260972 458798
rect 261220 443972 261248 468862
rect 261496 448526 261524 485046
rect 261588 468926 261616 485046
rect 261576 468920 261628 468926
rect 261576 468862 261628 468868
rect 281000 449478 281028 596702
rect 281552 487966 281580 700266
rect 283852 699825 283880 703520
rect 298836 700460 298888 700466
rect 298836 700402 298888 700408
rect 290556 700392 290608 700398
rect 290556 700334 290608 700340
rect 283838 699816 283894 699825
rect 283838 699751 283894 699760
rect 290464 696992 290516 696998
rect 290464 696934 290516 696940
rect 282368 597576 282420 597582
rect 282368 597518 282420 597524
rect 281632 597440 281684 597446
rect 281632 597382 281684 597388
rect 281644 596970 281672 597382
rect 281724 597304 281776 597310
rect 281724 597246 281776 597252
rect 281632 596964 281684 596970
rect 281632 596906 281684 596912
rect 281644 591394 281672 596906
rect 281736 596902 281764 597246
rect 282184 597236 282236 597242
rect 282184 597178 282236 597184
rect 282092 597168 282144 597174
rect 282092 597110 282144 597116
rect 281908 597032 281960 597038
rect 281908 596974 281960 596980
rect 281724 596896 281776 596902
rect 281724 596838 281776 596844
rect 281814 596864 281870 596873
rect 281632 591388 281684 591394
rect 281632 591330 281684 591336
rect 281632 591252 281684 591258
rect 281632 591194 281684 591200
rect 281540 487960 281592 487966
rect 281540 487902 281592 487908
rect 280988 449472 281040 449478
rect 280988 449414 281040 449420
rect 261484 448520 261536 448526
rect 261484 448462 261536 448468
rect 267096 448520 267148 448526
rect 267096 448462 267148 448468
rect 261496 443972 261524 448462
rect 265900 446888 265952 446894
rect 265900 446830 265952 446836
rect 264704 446820 264756 446826
rect 264704 446762 264756 446768
rect 264520 446752 264572 446758
rect 264520 446694 264572 446700
rect 261760 446412 261812 446418
rect 261760 446354 261812 446360
rect 261772 443972 261800 446354
rect 264426 446312 264482 446321
rect 264426 446247 264482 446256
rect 264242 444816 264298 444825
rect 264242 444751 264298 444760
rect 257436 443692 257488 443698
rect 257436 443634 257488 443640
rect 256976 443624 257028 443630
rect 256606 443592 256662 443601
rect 256542 443550 256606 443578
rect 256976 443566 257028 443572
rect 256606 443527 256662 443536
rect 256988 443494 257016 443566
rect 256976 443488 257028 443494
rect 257252 443488 257304 443494
rect 256976 443430 257028 443436
rect 257094 443436 257252 443442
rect 258906 443456 258962 443465
rect 257094 443430 257304 443436
rect 248880 443420 248932 443426
rect 243176 443362 243228 443368
rect 248880 443362 248932 443368
rect 248972 443420 249024 443426
rect 248972 443362 249024 443368
rect 249156 443420 249208 443426
rect 249366 443420 249576 443426
rect 249366 443414 249524 443420
rect 249156 443362 249208 443368
rect 249524 443362 249576 443368
rect 250812 443420 250864 443426
rect 250812 443362 250864 443368
rect 250904 443420 250956 443426
rect 250904 443362 250956 443368
rect 251732 443420 251784 443426
rect 257094 443414 257292 443430
rect 258750 443414 258906 443442
rect 259366 443456 259422 443465
rect 259302 443414 259366 443442
rect 258906 443391 258962 443400
rect 262126 443456 262182 443465
rect 262062 443414 262126 443442
rect 259366 443391 259422 443400
rect 262126 443391 262182 443400
rect 251732 443362 251784 443368
rect 203892 443352 203944 443358
rect 203720 443278 203826 443306
rect 203892 443294 203944 443300
rect 203720 441522 203748 443278
rect 263876 443080 263928 443086
rect 263876 443022 263928 443028
rect 263888 442474 263916 443022
rect 263876 442468 263928 442474
rect 263876 442410 263928 442416
rect 203708 441516 203760 441522
rect 203708 441458 203760 441464
rect 260010 400208 260066 400217
rect 260010 400143 260066 400152
rect 208214 398848 208270 398857
rect 208124 398812 208176 398818
rect 208214 398783 208270 398792
rect 208124 398754 208176 398760
rect 207940 398744 207992 398750
rect 207754 398712 207810 398721
rect 207940 398686 207992 398692
rect 207754 398647 207810 398656
rect 207664 398608 207716 398614
rect 206282 398576 206338 398585
rect 207664 398550 207716 398556
rect 206282 398511 206338 398520
rect 204994 397624 205050 397633
rect 204994 397559 205050 397568
rect 204904 395888 204956 395894
rect 204904 395830 204956 395836
rect 204260 351416 204312 351422
rect 204260 351358 204312 351364
rect 203616 215280 203668 215286
rect 203616 215222 203668 215228
rect 203524 33040 203576 33046
rect 203524 32982 203576 32988
rect 204272 16574 204300 351358
rect 203076 16546 203472 16574
rect 204272 16546 204852 16574
rect 202696 8016 202748 8022
rect 202696 7958 202748 7964
rect 202708 480 202736 7958
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 204824 3482 204852 16546
rect 204916 4010 204944 395830
rect 205008 355366 205036 397559
rect 205638 397080 205694 397089
rect 205638 397015 205694 397024
rect 204996 355360 205048 355366
rect 204996 355302 205048 355308
rect 205652 16574 205680 397015
rect 205652 16546 206232 16574
rect 204904 4004 204956 4010
rect 204904 3946 204956 3952
rect 204824 3454 205128 3482
rect 205100 480 205128 3454
rect 206204 480 206232 16546
rect 206296 4826 206324 398511
rect 207020 398472 207072 398478
rect 207020 398414 207072 398420
rect 206466 397488 206522 397497
rect 206466 397423 206522 397432
rect 206480 175982 206508 397423
rect 206468 175976 206520 175982
rect 206468 175918 206520 175924
rect 206284 4820 206336 4826
rect 206284 4762 206336 4768
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 398414
rect 207676 3670 207704 398550
rect 207664 3664 207716 3670
rect 207664 3606 207716 3612
rect 207768 3466 207796 398647
rect 207848 398540 207900 398546
rect 207848 398482 207900 398488
rect 207756 3460 207808 3466
rect 207756 3402 207808 3408
rect 207860 3398 207888 398482
rect 207952 5030 207980 398686
rect 208032 398676 208084 398682
rect 208032 398618 208084 398624
rect 208044 6322 208072 398618
rect 208136 37942 208164 398754
rect 208228 358086 208256 398783
rect 210238 398168 210294 398177
rect 210238 398103 210294 398112
rect 209780 398064 209832 398070
rect 209780 398006 209832 398012
rect 209136 397928 209188 397934
rect 209136 397870 209188 397876
rect 208398 394360 208454 394369
rect 208398 394295 208454 394304
rect 208216 358080 208268 358086
rect 208216 358022 208268 358028
rect 208124 37936 208176 37942
rect 208124 37878 208176 37884
rect 208412 16574 208440 394295
rect 209044 394256 209096 394262
rect 209044 394198 209096 394204
rect 208412 16546 208624 16574
rect 208032 6316 208084 6322
rect 208032 6258 208084 6264
rect 207940 5024 207992 5030
rect 207940 4966 207992 4972
rect 207848 3392 207900 3398
rect 207848 3334 207900 3340
rect 208596 480 208624 16546
rect 209056 3602 209084 394198
rect 209148 35222 209176 397870
rect 209228 397724 209280 397730
rect 209228 397666 209280 397672
rect 209240 171834 209268 397666
rect 209320 397520 209372 397526
rect 209320 397462 209372 397468
rect 209332 351218 209360 397462
rect 209792 396438 209820 398006
rect 210252 397633 210280 398103
rect 210344 397769 210372 400044
rect 210330 397760 210386 397769
rect 210330 397695 210386 397704
rect 210332 397656 210384 397662
rect 210238 397624 210294 397633
rect 210332 397598 210384 397604
rect 210238 397559 210294 397568
rect 210148 396772 210200 396778
rect 210148 396714 210200 396720
rect 209872 396704 209924 396710
rect 209872 396646 209924 396652
rect 209780 396432 209832 396438
rect 209780 396374 209832 396380
rect 209320 351212 209372 351218
rect 209320 351154 209372 351160
rect 209228 171828 209280 171834
rect 209228 171770 209280 171776
rect 209136 35216 209188 35222
rect 209136 35158 209188 35164
rect 209884 8974 209912 396646
rect 209964 396568 210016 396574
rect 209964 396510 210016 396516
rect 210056 396568 210108 396574
rect 210056 396510 210108 396516
rect 209976 9042 210004 396510
rect 210068 13190 210096 396510
rect 210056 13184 210108 13190
rect 210056 13126 210108 13132
rect 210160 13122 210188 396714
rect 210344 396386 210372 397598
rect 210436 396710 210464 400044
rect 210424 396704 210476 396710
rect 210424 396646 210476 396652
rect 210528 396642 210556 400044
rect 210620 396778 210648 400044
rect 210712 397984 210740 400044
rect 210804 398138 210832 400044
rect 210792 398132 210844 398138
rect 210792 398074 210844 398080
rect 210712 397956 210832 397984
rect 210698 397896 210754 397905
rect 210698 397831 210754 397840
rect 210608 396772 210660 396778
rect 210608 396714 210660 396720
rect 210516 396636 210568 396642
rect 210516 396578 210568 396584
rect 210608 396432 210660 396438
rect 210344 396358 210556 396386
rect 210608 396374 210660 396380
rect 210424 396092 210476 396098
rect 210424 396034 210476 396040
rect 210240 396024 210292 396030
rect 210240 395966 210292 395972
rect 210252 15910 210280 395966
rect 210240 15904 210292 15910
rect 210240 15846 210292 15852
rect 210148 13116 210200 13122
rect 210148 13058 210200 13064
rect 209964 9036 210016 9042
rect 209964 8978 210016 8984
rect 209872 8968 209924 8974
rect 209872 8910 209924 8916
rect 210436 4078 210464 396034
rect 210528 16046 210556 396358
rect 210620 177342 210648 396374
rect 210712 354006 210740 397831
rect 210804 397526 210832 397956
rect 210792 397520 210844 397526
rect 210792 397462 210844 397468
rect 210792 397384 210844 397390
rect 210792 397326 210844 397332
rect 210804 396098 210832 397326
rect 210792 396092 210844 396098
rect 210792 396034 210844 396040
rect 210896 393314 210924 400044
rect 210988 396574 211016 400044
rect 210976 396568 211028 396574
rect 210976 396510 211028 396516
rect 211080 396030 211108 400044
rect 211068 396024 211120 396030
rect 211068 395966 211120 395972
rect 211172 395321 211200 400044
rect 211264 397633 211292 400044
rect 211250 397624 211306 397633
rect 211250 397559 211306 397568
rect 211356 397497 211384 400044
rect 211448 397905 211476 400044
rect 211540 398449 211568 400044
rect 211526 398440 211582 398449
rect 211526 398375 211582 398384
rect 211434 397896 211490 397905
rect 211434 397831 211490 397840
rect 211632 397769 211660 400044
rect 211618 397760 211674 397769
rect 211618 397695 211674 397704
rect 211342 397488 211398 397497
rect 211342 397423 211398 397432
rect 211724 396794 211752 400044
rect 211252 396772 211304 396778
rect 211252 396714 211304 396720
rect 211540 396766 211752 396794
rect 211158 395312 211214 395321
rect 211158 395247 211214 395256
rect 210804 393286 210924 393314
rect 210700 354000 210752 354006
rect 210700 353942 210752 353948
rect 210608 177336 210660 177342
rect 210608 177278 210660 177284
rect 210516 16040 210568 16046
rect 210516 15982 210568 15988
rect 210804 9110 210832 393286
rect 211264 11762 211292 396714
rect 211344 396636 211396 396642
rect 211344 396578 211396 396584
rect 211356 14550 211384 396578
rect 211436 396568 211488 396574
rect 211436 396510 211488 396516
rect 211448 14618 211476 396510
rect 211436 14612 211488 14618
rect 211436 14554 211488 14560
rect 211344 14544 211396 14550
rect 211344 14486 211396 14492
rect 211540 14482 211568 396766
rect 211620 396704 211672 396710
rect 211816 396658 211844 400044
rect 211908 396710 211936 400044
rect 212000 396778 212028 400044
rect 211988 396772 212040 396778
rect 211988 396714 212040 396720
rect 211620 396646 211672 396652
rect 211632 354142 211660 396646
rect 211724 396630 211844 396658
rect 211896 396704 211948 396710
rect 211896 396646 211948 396652
rect 212092 396642 212120 400044
rect 212184 398857 212212 400044
rect 212170 398848 212226 398857
rect 212170 398783 212226 398792
rect 212172 398744 212224 398750
rect 212172 398686 212224 398692
rect 212184 398002 212212 398686
rect 212276 398410 212304 400044
rect 212264 398404 212316 398410
rect 212264 398346 212316 398352
rect 212172 397996 212224 398002
rect 212172 397938 212224 397944
rect 212262 397760 212318 397769
rect 212262 397695 212318 397704
rect 212172 397520 212224 397526
rect 212172 397462 212224 397468
rect 212080 396636 212132 396642
rect 211620 354136 211672 354142
rect 211620 354078 211672 354084
rect 211724 354074 211752 396630
rect 212080 396578 212132 396584
rect 212184 396522 212212 397462
rect 211816 396494 212212 396522
rect 211712 354068 211764 354074
rect 211712 354010 211764 354016
rect 211620 46300 211672 46306
rect 211620 46242 211672 46248
rect 211632 16574 211660 46242
rect 211632 16546 211752 16574
rect 211528 14476 211580 14482
rect 211528 14418 211580 14424
rect 211252 11756 211304 11762
rect 211252 11698 211304 11704
rect 210792 9104 210844 9110
rect 210792 9046 210844 9052
rect 210976 4820 211028 4826
rect 210976 4762 211028 4768
rect 210424 4072 210476 4078
rect 210424 4014 210476 4020
rect 209044 3596 209096 3602
rect 209044 3538 209096 3544
rect 209780 3596 209832 3602
rect 209780 3538 209832 3544
rect 209792 480 209820 3538
rect 210988 480 211016 4762
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 14686 211844 396494
rect 212276 393314 212304 397695
rect 211908 393286 212304 393314
rect 211908 354346 211936 393286
rect 211896 354340 211948 354346
rect 211896 354282 211948 354288
rect 211804 14680 211856 14686
rect 211804 14622 211856 14628
rect 212368 11830 212396 400044
rect 212460 396574 212488 400044
rect 212552 397497 212580 400044
rect 212644 398721 212672 400044
rect 212630 398712 212686 398721
rect 212630 398647 212686 398656
rect 212632 398404 212684 398410
rect 212632 398346 212684 398352
rect 212644 398070 212672 398346
rect 212632 398064 212684 398070
rect 212632 398006 212684 398012
rect 212630 397896 212686 397905
rect 212630 397831 212686 397840
rect 212538 397488 212594 397497
rect 212538 397423 212594 397432
rect 212540 397248 212592 397254
rect 212540 397190 212592 397196
rect 212552 396846 212580 397190
rect 212540 396840 212592 396846
rect 212540 396782 212592 396788
rect 212448 396568 212500 396574
rect 212448 396510 212500 396516
rect 212644 396386 212672 397831
rect 212736 397497 212764 400044
rect 212828 398585 212856 400044
rect 212814 398576 212870 398585
rect 212814 398511 212870 398520
rect 212920 397594 212948 400044
rect 212908 397588 212960 397594
rect 212908 397530 212960 397536
rect 212722 397488 212778 397497
rect 212722 397423 212778 397432
rect 212908 397452 212960 397458
rect 212908 397394 212960 397400
rect 212920 397050 212948 397394
rect 213012 397050 213040 400044
rect 212908 397044 212960 397050
rect 212908 396986 212960 396992
rect 213000 397044 213052 397050
rect 213000 396986 213052 396992
rect 213104 396794 213132 400044
rect 212724 396772 212776 396778
rect 212724 396714 212776 396720
rect 212828 396766 213132 396794
rect 212460 396358 212672 396386
rect 212460 393990 212488 396358
rect 212448 393984 212500 393990
rect 212448 393926 212500 393932
rect 212736 12034 212764 396714
rect 212828 15978 212856 396766
rect 213000 396704 213052 396710
rect 213196 396658 213224 400044
rect 213288 397322 213316 400044
rect 213380 398041 213408 400044
rect 213366 398032 213422 398041
rect 213366 397967 213422 397976
rect 213472 397712 213500 400044
rect 213380 397684 213500 397712
rect 213276 397316 213328 397322
rect 213276 397258 213328 397264
rect 213380 397254 213408 397684
rect 213460 397588 213512 397594
rect 213460 397530 213512 397536
rect 213368 397248 213420 397254
rect 213368 397190 213420 397196
rect 213368 397044 213420 397050
rect 213368 396986 213420 396992
rect 213000 396646 213052 396652
rect 212908 396636 212960 396642
rect 212908 396578 212960 396584
rect 212920 354210 212948 396578
rect 213012 354278 213040 396646
rect 213104 396630 213224 396658
rect 213000 354272 213052 354278
rect 213000 354214 213052 354220
rect 212908 354204 212960 354210
rect 212908 354146 212960 354152
rect 212816 15972 212868 15978
rect 212816 15914 212868 15920
rect 212724 12028 212776 12034
rect 212724 11970 212776 11976
rect 213104 11966 213132 396630
rect 213184 396432 213236 396438
rect 213184 396374 213236 396380
rect 213092 11960 213144 11966
rect 213092 11902 213144 11908
rect 212356 11824 212408 11830
rect 212356 11766 212408 11772
rect 213196 3806 213224 396374
rect 213276 394936 213328 394942
rect 213276 394878 213328 394884
rect 213288 355502 213316 394878
rect 213380 392630 213408 396986
rect 213368 392624 213420 392630
rect 213368 392566 213420 392572
rect 213276 355496 213328 355502
rect 213276 355438 213328 355444
rect 213276 352572 213328 352578
rect 213276 352514 213328 352520
rect 213184 3800 213236 3806
rect 213184 3742 213236 3748
rect 213288 3602 213316 352514
rect 213472 11898 213500 397530
rect 213564 396642 213592 400044
rect 213656 396710 213684 400044
rect 213748 396778 213776 400044
rect 213840 397526 213868 400044
rect 213932 398177 213960 400044
rect 213918 398168 213974 398177
rect 213918 398103 213974 398112
rect 214024 397905 214052 400044
rect 214010 397896 214066 397905
rect 214010 397831 214066 397840
rect 213920 397588 213972 397594
rect 213920 397530 213972 397536
rect 213828 397520 213880 397526
rect 213828 397462 213880 397468
rect 213932 397338 213960 397530
rect 214116 397474 214144 400044
rect 214208 397497 214236 400044
rect 214300 397633 214328 400044
rect 214286 397624 214342 397633
rect 214286 397559 214342 397568
rect 213840 397310 213960 397338
rect 214024 397446 214144 397474
rect 214194 397488 214250 397497
rect 213736 396772 213788 396778
rect 213736 396714 213788 396720
rect 213644 396704 213696 396710
rect 213644 396646 213696 396652
rect 213552 396636 213604 396642
rect 213552 396578 213604 396584
rect 213840 394942 213868 397310
rect 214024 396681 214052 397446
rect 214194 397423 214250 397432
rect 214104 397044 214156 397050
rect 214104 396986 214156 396992
rect 214010 396672 214066 396681
rect 214010 396607 214066 396616
rect 213920 396500 213972 396506
rect 213920 396442 213972 396448
rect 213828 394936 213880 394942
rect 213828 394878 213880 394884
rect 213460 11892 213512 11898
rect 213460 11834 213512 11840
rect 213932 4962 213960 396442
rect 214012 395004 214064 395010
rect 214012 394946 214064 394952
rect 213920 4956 213972 4962
rect 213920 4898 213972 4904
rect 214024 4894 214052 394946
rect 214116 9178 214144 396986
rect 214392 396658 214420 400044
rect 214196 396636 214248 396642
rect 214196 396578 214248 396584
rect 214300 396630 214420 396658
rect 214208 9246 214236 396578
rect 214300 13258 214328 396630
rect 214380 396568 214432 396574
rect 214380 396510 214432 396516
rect 214392 13462 214420 396510
rect 214484 395622 214512 400044
rect 214576 397050 214604 400044
rect 214564 397044 214616 397050
rect 214564 396986 214616 396992
rect 214668 396658 214696 400044
rect 214760 397769 214788 400044
rect 214746 397760 214802 397769
rect 214746 397695 214802 397704
rect 214746 397624 214802 397633
rect 214746 397559 214802 397568
rect 214576 396630 214696 396658
rect 214472 395616 214524 395622
rect 214472 395558 214524 395564
rect 214472 395480 214524 395486
rect 214472 395422 214524 395428
rect 214380 13456 214432 13462
rect 214380 13398 214432 13404
rect 214484 13394 214512 395422
rect 214472 13388 214524 13394
rect 214472 13330 214524 13336
rect 214576 13326 214604 396630
rect 214656 395616 214708 395622
rect 214656 395558 214708 395564
rect 214668 352646 214696 395558
rect 214760 395418 214788 397559
rect 214748 395412 214800 395418
rect 214748 395354 214800 395360
rect 214852 395010 214880 400044
rect 214944 395486 214972 400044
rect 215036 396506 215064 400044
rect 215128 396642 215156 400044
rect 215116 396636 215168 396642
rect 215116 396578 215168 396584
rect 215220 396574 215248 400044
rect 215312 398041 215340 400044
rect 215298 398032 215354 398041
rect 215298 397967 215354 397976
rect 215300 397860 215352 397866
rect 215300 397802 215352 397808
rect 215312 397118 215340 397802
rect 215404 397497 215432 400044
rect 215496 397633 215524 400044
rect 215588 397769 215616 400044
rect 215574 397760 215630 397769
rect 215574 397695 215630 397704
rect 215482 397624 215538 397633
rect 215482 397559 215538 397568
rect 215390 397488 215446 397497
rect 215390 397423 215446 397432
rect 215300 397112 215352 397118
rect 215300 397054 215352 397060
rect 215680 396930 215708 400044
rect 215772 397497 215800 400044
rect 215864 397662 215892 400044
rect 215852 397656 215904 397662
rect 215852 397598 215904 397604
rect 215758 397488 215814 397497
rect 215758 397423 215814 397432
rect 215404 396902 215708 396930
rect 215300 396840 215352 396846
rect 215300 396782 215352 396788
rect 215208 396568 215260 396574
rect 215208 396510 215260 396516
rect 215024 396500 215076 396506
rect 215024 396442 215076 396448
rect 215312 396438 215340 396782
rect 215300 396432 215352 396438
rect 215300 396374 215352 396380
rect 214932 395480 214984 395486
rect 214932 395422 214984 395428
rect 214840 395004 214892 395010
rect 214840 394946 214892 394952
rect 214656 352640 214708 352646
rect 214656 352582 214708 352588
rect 214564 13320 214616 13326
rect 214564 13262 214616 13268
rect 214288 13252 214340 13258
rect 214288 13194 214340 13200
rect 215404 10334 215432 396902
rect 215956 396778 215984 400044
rect 215484 396772 215536 396778
rect 215484 396714 215536 396720
rect 215944 396772 215996 396778
rect 215944 396714 215996 396720
rect 215496 10402 215524 396714
rect 216048 396658 216076 400044
rect 215760 396636 215812 396642
rect 215760 396578 215812 396584
rect 215864 396630 216076 396658
rect 215576 396568 215628 396574
rect 215576 396510 215628 396516
rect 215588 13530 215616 396510
rect 215668 396364 215720 396370
rect 215668 396306 215720 396312
rect 215680 14754 215708 396306
rect 215772 354414 215800 396578
rect 215864 355434 215892 396630
rect 216140 396370 216168 400044
rect 216128 396364 216180 396370
rect 216128 396306 216180 396312
rect 216232 396250 216260 400044
rect 216324 398154 216352 400044
rect 216416 398410 216444 400044
rect 216404 398404 216456 398410
rect 216404 398346 216456 398352
rect 216324 398126 216444 398154
rect 216312 398064 216364 398070
rect 216312 398006 216364 398012
rect 216140 396222 216260 396250
rect 215944 395684 215996 395690
rect 215944 395626 215996 395632
rect 215956 392698 215984 395626
rect 215944 392692 215996 392698
rect 215944 392634 215996 392640
rect 215852 355428 215904 355434
rect 215852 355370 215904 355376
rect 215760 354408 215812 354414
rect 215760 354350 215812 354356
rect 215760 177336 215812 177342
rect 215760 177278 215812 177284
rect 215668 14748 215720 14754
rect 215668 14690 215720 14696
rect 215576 13524 215628 13530
rect 215576 13466 215628 13472
rect 215484 10396 215536 10402
rect 215484 10338 215536 10344
rect 215392 10328 215444 10334
rect 215392 10270 215444 10276
rect 214196 9240 214248 9246
rect 214196 9182 214248 9188
rect 214104 9172 214156 9178
rect 214104 9114 214156 9120
rect 215772 6914 215800 177278
rect 216140 10470 216168 396222
rect 216324 395690 216352 398006
rect 216312 395684 216364 395690
rect 216312 395626 216364 395632
rect 216416 395350 216444 398126
rect 216508 396642 216536 400044
rect 216496 396636 216548 396642
rect 216496 396578 216548 396584
rect 216600 396574 216628 400044
rect 216692 397769 216720 400044
rect 216784 398993 216812 400044
rect 216770 398984 216826 398993
rect 216770 398919 216826 398928
rect 216772 398880 216824 398886
rect 216772 398822 216824 398828
rect 216678 397760 216734 397769
rect 216678 397695 216734 397704
rect 216784 396794 216812 398822
rect 216876 397633 216904 400044
rect 216862 397624 216918 397633
rect 216862 397559 216918 397568
rect 216968 397497 216996 400044
rect 216954 397488 217010 397497
rect 216954 397423 217010 397432
rect 216692 396766 216812 396794
rect 216588 396568 216640 396574
rect 216588 396510 216640 396516
rect 216692 395554 216720 396766
rect 217060 396658 217088 400044
rect 217152 397905 217180 400044
rect 217138 397896 217194 397905
rect 217138 397831 217194 397840
rect 217244 397594 217272 400044
rect 217232 397588 217284 397594
rect 217232 397530 217284 397536
rect 216784 396630 217088 396658
rect 216680 395548 216732 395554
rect 216680 395490 216732 395496
rect 216404 395344 216456 395350
rect 216404 395286 216456 395292
rect 216784 10538 216812 396630
rect 216864 396568 216916 396574
rect 217336 396522 217364 400044
rect 216864 396510 216916 396516
rect 216876 10742 216904 396510
rect 216968 396494 217364 396522
rect 216864 10736 216916 10742
rect 216864 10678 216916 10684
rect 216968 10606 216996 396494
rect 217048 396432 217100 396438
rect 217048 396374 217100 396380
rect 217060 10674 217088 396374
rect 217232 396364 217284 396370
rect 217232 396306 217284 396312
rect 217140 396296 217192 396302
rect 217140 396238 217192 396244
rect 217152 14822 217180 396238
rect 217244 14890 217272 396306
rect 217428 396302 217456 400044
rect 217416 396296 217468 396302
rect 217416 396238 217468 396244
rect 217520 396114 217548 400044
rect 217612 396438 217640 400044
rect 217704 398886 217732 400044
rect 217692 398880 217744 398886
rect 217692 398822 217744 398828
rect 217692 398676 217744 398682
rect 217692 398618 217744 398624
rect 217600 396432 217652 396438
rect 217600 396374 217652 396380
rect 217520 396086 217640 396114
rect 217324 396024 217376 396030
rect 217324 395966 217376 395972
rect 217232 14884 217284 14890
rect 217232 14826 217284 14832
rect 217140 14816 217192 14822
rect 217140 14758 217192 14764
rect 217048 10668 217100 10674
rect 217048 10610 217100 10616
rect 216956 10600 217008 10606
rect 216956 10542 217008 10548
rect 216772 10532 216824 10538
rect 216772 10474 216824 10480
rect 216128 10464 216180 10470
rect 216128 10406 216180 10412
rect 217336 7614 217364 395966
rect 217612 393394 217640 396086
rect 217704 396030 217732 398618
rect 217796 397934 217824 400044
rect 217784 397928 217836 397934
rect 217784 397870 217836 397876
rect 217888 396574 217916 400044
rect 217876 396568 217928 396574
rect 217876 396510 217928 396516
rect 217980 396370 218008 400044
rect 218072 397769 218100 400044
rect 218058 397760 218114 397769
rect 218058 397695 218114 397704
rect 218164 397497 218192 400044
rect 218256 397633 218284 400044
rect 218348 397730 218376 400044
rect 218336 397724 218388 397730
rect 218336 397666 218388 397672
rect 218242 397624 218298 397633
rect 218242 397559 218298 397568
rect 218150 397488 218206 397497
rect 218150 397423 218206 397432
rect 218060 397044 218112 397050
rect 218060 396986 218112 396992
rect 217968 396364 218020 396370
rect 217968 396306 218020 396312
rect 217692 396024 217744 396030
rect 217692 395966 217744 395972
rect 218072 395826 218100 396986
rect 218440 396930 218468 400044
rect 218152 396908 218204 396914
rect 218152 396850 218204 396856
rect 218348 396902 218468 396930
rect 218060 395820 218112 395826
rect 218060 395762 218112 395768
rect 218164 395758 218192 396850
rect 218244 396636 218296 396642
rect 218244 396578 218296 396584
rect 218152 395752 218204 395758
rect 218152 395694 218204 395700
rect 217520 393366 217640 393394
rect 217324 7608 217376 7614
rect 217324 7550 217376 7556
rect 215680 6886 215800 6914
rect 214012 4888 214064 4894
rect 214012 4830 214064 4836
rect 214472 4888 214524 4894
rect 214472 4830 214524 4836
rect 213276 3596 213328 3602
rect 213276 3538 213328 3544
rect 213368 3052 213420 3058
rect 213368 2994 213420 3000
rect 213380 480 213408 2994
rect 214484 480 214512 4830
rect 215680 480 215708 6886
rect 217520 6254 217548 393366
rect 218256 12238 218284 396578
rect 218348 396574 218376 396902
rect 218428 396772 218480 396778
rect 218428 396714 218480 396720
rect 218336 396568 218388 396574
rect 218336 396510 218388 396516
rect 218336 396364 218388 396370
rect 218336 396306 218388 396312
rect 218244 12232 218296 12238
rect 218244 12174 218296 12180
rect 218348 12170 218376 396306
rect 218440 15026 218468 396714
rect 218532 396658 218560 400044
rect 218624 396778 218652 400044
rect 218612 396772 218664 396778
rect 218612 396714 218664 396720
rect 218716 396658 218744 400044
rect 218808 396914 218836 400044
rect 218900 398002 218928 400044
rect 218888 397996 218940 398002
rect 218888 397938 218940 397944
rect 218886 397896 218942 397905
rect 218886 397831 218942 397840
rect 218900 397050 218928 397831
rect 218888 397044 218940 397050
rect 218888 396986 218940 396992
rect 218796 396908 218848 396914
rect 218796 396850 218848 396856
rect 218532 396630 218652 396658
rect 218716 396630 218928 396658
rect 218520 396432 218572 396438
rect 218520 396374 218572 396380
rect 218428 15020 218480 15026
rect 218428 14962 218480 14968
rect 218532 14958 218560 396374
rect 218624 352714 218652 396630
rect 218796 396568 218848 396574
rect 218796 396510 218848 396516
rect 218704 396500 218756 396506
rect 218704 396442 218756 396448
rect 218716 355570 218744 396442
rect 218704 355564 218756 355570
rect 218704 355506 218756 355512
rect 218612 352708 218664 352714
rect 218612 352650 218664 352656
rect 218520 14952 218572 14958
rect 218520 14894 218572 14900
rect 218336 12164 218388 12170
rect 218336 12106 218388 12112
rect 218808 10810 218836 396510
rect 218900 12102 218928 396630
rect 218992 396370 219020 400044
rect 219084 396438 219112 400044
rect 219176 396506 219204 400044
rect 219268 396642 219296 400044
rect 219360 398449 219388 400044
rect 219452 398750 219480 400044
rect 219440 398744 219492 398750
rect 219440 398686 219492 398692
rect 219346 398440 219402 398449
rect 219346 398375 219402 398384
rect 219346 398304 219402 398313
rect 219346 398239 219402 398248
rect 219256 396636 219308 396642
rect 219256 396578 219308 396584
rect 219164 396500 219216 396506
rect 219164 396442 219216 396448
rect 219072 396432 219124 396438
rect 219072 396374 219124 396380
rect 218980 396364 219032 396370
rect 218980 396306 219032 396312
rect 219360 395865 219388 398239
rect 219544 397633 219572 400044
rect 219636 397769 219664 400044
rect 219728 398682 219756 400044
rect 219716 398676 219768 398682
rect 219716 398618 219768 398624
rect 219820 398313 219848 400044
rect 219806 398304 219862 398313
rect 219806 398239 219862 398248
rect 219622 397760 219678 397769
rect 219622 397695 219678 397704
rect 219624 397656 219676 397662
rect 219530 397624 219586 397633
rect 219624 397598 219676 397604
rect 219530 397559 219586 397568
rect 219440 396908 219492 396914
rect 219440 396850 219492 396856
rect 219346 395856 219402 395865
rect 219346 395791 219402 395800
rect 219452 394262 219480 396850
rect 219636 396692 219664 397598
rect 219912 397497 219940 400044
rect 220004 398818 220032 400044
rect 219992 398812 220044 398818
rect 219992 398754 220044 398760
rect 219992 397724 220044 397730
rect 219992 397666 220044 397672
rect 219898 397488 219954 397497
rect 219898 397423 219954 397432
rect 219716 396840 219768 396846
rect 219716 396782 219768 396788
rect 219544 396664 219664 396692
rect 219440 394256 219492 394262
rect 219440 394198 219492 394204
rect 219440 393984 219492 393990
rect 219440 393926 219492 393932
rect 218888 12096 218940 12102
rect 218888 12038 218940 12044
rect 218796 10804 218848 10810
rect 218796 10746 218848 10752
rect 217508 6248 217560 6254
rect 217508 6190 217560 6196
rect 219256 4072 219308 4078
rect 219256 4014 219308 4020
rect 218060 3868 218112 3874
rect 218060 3810 218112 3816
rect 216864 3664 216916 3670
rect 216864 3606 216916 3612
rect 216876 480 216904 3606
rect 218072 480 218100 3810
rect 219268 480 219296 4014
rect 219452 490 219480 393926
rect 219544 3534 219572 396664
rect 219624 396568 219676 396574
rect 219624 396510 219676 396516
rect 219636 5370 219664 396510
rect 219624 5364 219676 5370
rect 219624 5306 219676 5312
rect 219728 5098 219756 396782
rect 219808 396636 219860 396642
rect 219808 396578 219860 396584
rect 219820 6390 219848 396578
rect 219900 396500 219952 396506
rect 219900 396442 219952 396448
rect 219912 177410 219940 396442
rect 220004 396352 220032 397666
rect 220096 396914 220124 400044
rect 220084 396908 220136 396914
rect 220084 396850 220136 396856
rect 220188 396846 220216 400044
rect 220176 396840 220228 396846
rect 220176 396782 220228 396788
rect 220280 396506 220308 400044
rect 220372 397662 220400 400044
rect 220360 397656 220412 397662
rect 220360 397598 220412 397604
rect 220360 397520 220412 397526
rect 220360 397462 220412 397468
rect 220268 396500 220320 396506
rect 220268 396442 220320 396448
rect 220004 396324 220216 396352
rect 219992 396228 220044 396234
rect 219992 396170 220044 396176
rect 220004 177478 220032 396170
rect 220084 396024 220136 396030
rect 220084 395966 220136 395972
rect 219992 177472 220044 177478
rect 219992 177414 220044 177420
rect 219900 177404 219952 177410
rect 219900 177346 219952 177352
rect 219808 6384 219860 6390
rect 219808 6326 219860 6332
rect 219716 5092 219768 5098
rect 219716 5034 219768 5040
rect 219532 3528 219584 3534
rect 219532 3470 219584 3476
rect 220096 3058 220124 395966
rect 220188 393990 220216 396324
rect 220176 393984 220228 393990
rect 220176 393926 220228 393932
rect 220372 393314 220400 397462
rect 220464 396642 220492 400044
rect 220556 396710 220584 400044
rect 220544 396704 220596 396710
rect 220544 396646 220596 396652
rect 220452 396636 220504 396642
rect 220452 396578 220504 396584
rect 220648 396574 220676 400044
rect 220636 396568 220688 396574
rect 220636 396510 220688 396516
rect 220740 396234 220768 400044
rect 220832 397769 220860 400044
rect 220818 397760 220874 397769
rect 220818 397695 220874 397704
rect 220820 397656 220872 397662
rect 220820 397598 220872 397604
rect 220728 396228 220780 396234
rect 220728 396170 220780 396176
rect 220188 393286 220400 393314
rect 220188 16114 220216 393286
rect 220176 16108 220228 16114
rect 220176 16050 220228 16056
rect 220832 4078 220860 397598
rect 220924 397526 220952 400044
rect 220912 397520 220964 397526
rect 221016 397497 221044 400044
rect 220912 397462 220964 397468
rect 221002 397488 221058 397497
rect 221002 397423 221058 397432
rect 221108 396817 221136 400044
rect 221200 398138 221228 400044
rect 221188 398132 221240 398138
rect 221188 398074 221240 398080
rect 221292 397633 221320 400044
rect 221278 397624 221334 397633
rect 221278 397559 221334 397568
rect 221094 396808 221150 396817
rect 221094 396743 221150 396752
rect 221096 396704 221148 396710
rect 221384 396692 221412 400044
rect 221096 396646 221148 396652
rect 221200 396664 221412 396692
rect 221004 396636 221056 396642
rect 221004 396578 221056 396584
rect 220912 396228 220964 396234
rect 220912 396170 220964 396176
rect 220924 5234 220952 396170
rect 221016 7750 221044 396578
rect 221004 7744 221056 7750
rect 221004 7686 221056 7692
rect 221108 7682 221136 396646
rect 221200 9314 221228 396664
rect 221280 396568 221332 396574
rect 221280 396510 221332 396516
rect 221292 9382 221320 396510
rect 221372 396500 221424 396506
rect 221372 396442 221424 396448
rect 221384 351286 221412 396442
rect 221476 394058 221504 400044
rect 221568 396710 221596 400044
rect 221660 396982 221688 400044
rect 221648 396976 221700 396982
rect 221648 396918 221700 396924
rect 221556 396704 221608 396710
rect 221556 396646 221608 396652
rect 221464 394052 221516 394058
rect 221464 393994 221516 394000
rect 221752 393314 221780 400044
rect 221844 396642 221872 400044
rect 221832 396636 221884 396642
rect 221832 396578 221884 396584
rect 221936 396574 221964 400044
rect 221924 396568 221976 396574
rect 221924 396510 221976 396516
rect 222028 396234 222056 400044
rect 222120 396506 222148 400044
rect 222212 397594 222240 400044
rect 222200 397588 222252 397594
rect 222200 397530 222252 397536
rect 222304 397497 222332 400044
rect 222396 397633 222424 400044
rect 222382 397624 222438 397633
rect 222382 397559 222438 397568
rect 222384 397520 222436 397526
rect 222290 397488 222346 397497
rect 222384 397462 222436 397468
rect 222290 397423 222346 397432
rect 222396 397066 222424 397462
rect 222304 397038 222424 397066
rect 222108 396500 222160 396506
rect 222108 396442 222160 396448
rect 222016 396228 222068 396234
rect 222016 396170 222068 396176
rect 221568 393286 221780 393314
rect 221372 351280 221424 351286
rect 221372 351222 221424 351228
rect 221280 9376 221332 9382
rect 221280 9318 221332 9324
rect 221188 9308 221240 9314
rect 221188 9250 221240 9256
rect 221096 7676 221148 7682
rect 221096 7618 221148 7624
rect 220912 5228 220964 5234
rect 220912 5170 220964 5176
rect 221568 5166 221596 393286
rect 221556 5160 221608 5166
rect 221556 5102 221608 5108
rect 220820 4072 220872 4078
rect 220820 4014 220872 4020
rect 222304 3670 222332 397038
rect 222384 396908 222436 396914
rect 222384 396850 222436 396856
rect 222396 7818 222424 396850
rect 222488 396692 222516 400044
rect 222580 396846 222608 400044
rect 222672 396914 222700 400044
rect 222660 396908 222712 396914
rect 222660 396850 222712 396856
rect 222568 396840 222620 396846
rect 222764 396794 222792 400044
rect 222856 398614 222884 400044
rect 222844 398608 222896 398614
rect 222844 398550 222896 398556
rect 222568 396782 222620 396788
rect 222672 396766 222792 396794
rect 222844 396840 222896 396846
rect 222844 396782 222896 396788
rect 222488 396664 222608 396692
rect 222476 396568 222528 396574
rect 222476 396510 222528 396516
rect 222488 7886 222516 396510
rect 222580 9450 222608 396664
rect 222672 46238 222700 396766
rect 222856 393314 222884 396782
rect 222764 393286 222884 393314
rect 222764 352782 222792 393286
rect 222752 352776 222804 352782
rect 222752 352718 222804 352724
rect 222752 350600 222804 350606
rect 222752 350542 222804 350548
rect 222660 46232 222712 46238
rect 222660 46174 222712 46180
rect 222568 9444 222620 9450
rect 222568 9386 222620 9392
rect 222476 7880 222528 7886
rect 222476 7822 222528 7828
rect 222384 7812 222436 7818
rect 222384 7754 222436 7760
rect 222292 3664 222344 3670
rect 222292 3606 222344 3612
rect 220084 3052 220136 3058
rect 220084 2994 220136 3000
rect 221556 3052 221608 3058
rect 221556 2994 221608 3000
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 219452 462 220032 490
rect 221568 480 221596 2994
rect 222764 480 222792 350542
rect 222948 5302 222976 400044
rect 223040 397866 223068 400044
rect 223132 398070 223160 400044
rect 223120 398064 223172 398070
rect 223120 398006 223172 398012
rect 223028 397860 223080 397866
rect 223028 397802 223080 397808
rect 223224 393314 223252 400044
rect 223316 396574 223344 400044
rect 223408 396778 223436 400044
rect 223396 396772 223448 396778
rect 223396 396714 223448 396720
rect 223304 396568 223356 396574
rect 223304 396510 223356 396516
rect 223500 394126 223528 400044
rect 223592 397633 223620 400044
rect 223684 398274 223712 400044
rect 223672 398268 223724 398274
rect 223672 398210 223724 398216
rect 223776 397905 223804 400044
rect 223762 397896 223818 397905
rect 223762 397831 223818 397840
rect 223578 397624 223634 397633
rect 223578 397559 223634 397568
rect 223868 397497 223896 400044
rect 223960 397769 223988 400044
rect 223946 397760 224002 397769
rect 223946 397695 224002 397704
rect 223854 397488 223910 397497
rect 223854 397423 223910 397432
rect 223856 396840 223908 396846
rect 223856 396782 223908 396788
rect 223764 396636 223816 396642
rect 223764 396578 223816 396584
rect 223488 394120 223540 394126
rect 223488 394062 223540 394068
rect 223224 393286 223528 393314
rect 223500 5438 223528 393286
rect 223776 6662 223804 396578
rect 223764 6656 223816 6662
rect 223764 6598 223816 6604
rect 223868 6526 223896 396782
rect 224052 396692 224080 400044
rect 223960 396664 224080 396692
rect 223856 6520 223908 6526
rect 223856 6462 223908 6468
rect 223960 6458 223988 396664
rect 224040 396568 224092 396574
rect 224040 396510 224092 396516
rect 224052 17270 224080 396510
rect 224144 395894 224172 400044
rect 224132 395888 224184 395894
rect 224132 395830 224184 395836
rect 224132 394188 224184 394194
rect 224132 394130 224184 394136
rect 224144 351354 224172 394130
rect 224132 351348 224184 351354
rect 224132 351290 224184 351296
rect 224040 17264 224092 17270
rect 224040 17206 224092 17212
rect 223948 6452 224000 6458
rect 223948 6394 224000 6400
rect 223488 5432 223540 5438
rect 223488 5374 223540 5380
rect 222936 5296 222988 5302
rect 222936 5238 222988 5244
rect 224236 3738 224264 400044
rect 224328 396846 224356 400044
rect 224316 396840 224368 396846
rect 224316 396782 224368 396788
rect 224316 396704 224368 396710
rect 224316 396646 224368 396652
rect 224328 391270 224356 396646
rect 224420 396574 224448 400044
rect 224408 396568 224460 396574
rect 224408 396510 224460 396516
rect 224512 394194 224540 400044
rect 224500 394188 224552 394194
rect 224500 394130 224552 394136
rect 224604 393314 224632 400044
rect 224696 397390 224724 400044
rect 224684 397384 224736 397390
rect 224684 397326 224736 397332
rect 224788 396710 224816 400044
rect 224776 396704 224828 396710
rect 224776 396646 224828 396652
rect 224880 396642 224908 400044
rect 224972 397633 225000 400044
rect 225064 398342 225092 400044
rect 225156 398546 225184 400044
rect 225144 398540 225196 398546
rect 225144 398482 225196 398488
rect 225052 398336 225104 398342
rect 225052 398278 225104 398284
rect 224958 397624 225014 397633
rect 224958 397559 225014 397568
rect 225248 396953 225276 400044
rect 225234 396944 225290 396953
rect 225234 396879 225290 396888
rect 224868 396636 224920 396642
rect 224868 396578 224920 396584
rect 225340 394074 225368 400044
rect 225432 397497 225460 400044
rect 225418 397488 225474 397497
rect 225418 397423 225474 397432
rect 224420 393286 224632 393314
rect 225064 394046 225368 394074
rect 224316 391264 224368 391270
rect 224316 391206 224368 391212
rect 224420 6594 224448 393286
rect 224408 6588 224460 6594
rect 224408 6530 224460 6536
rect 225064 3942 225092 394046
rect 225524 393972 225552 400044
rect 225616 394262 225644 400044
rect 225604 394256 225656 394262
rect 225604 394198 225656 394204
rect 225340 393944 225552 393972
rect 225604 393984 225656 393990
rect 225144 393916 225196 393922
rect 225144 393858 225196 393864
rect 225156 6186 225184 393858
rect 225236 393780 225288 393786
rect 225236 393722 225288 393728
rect 225248 8022 225276 393722
rect 225236 8016 225288 8022
rect 225236 7958 225288 7964
rect 225340 7954 225368 393944
rect 225604 393926 225656 393932
rect 225512 393848 225564 393854
rect 225512 393790 225564 393796
rect 225420 391740 225472 391746
rect 225420 391682 225472 391688
rect 225432 177546 225460 391682
rect 225524 177614 225552 393790
rect 225616 351422 225644 393926
rect 225708 393922 225736 400044
rect 225800 397186 225828 400044
rect 225788 397180 225840 397186
rect 225788 397122 225840 397128
rect 225696 393916 225748 393922
rect 225696 393858 225748 393864
rect 225892 389174 225920 400044
rect 225984 391746 226012 400044
rect 226076 393786 226104 400044
rect 226168 393854 226196 400044
rect 226260 393990 226288 400044
rect 226352 397089 226380 400044
rect 226444 398478 226472 400044
rect 226432 398472 226484 398478
rect 226432 398414 226484 398420
rect 226432 397520 226484 397526
rect 226536 397497 226564 400044
rect 226432 397462 226484 397468
rect 226522 397488 226578 397497
rect 226338 397080 226394 397089
rect 226338 397015 226394 397024
rect 226444 394346 226472 397462
rect 226522 397423 226578 397432
rect 226352 394318 226472 394346
rect 226248 393984 226300 393990
rect 226248 393926 226300 393932
rect 226156 393848 226208 393854
rect 226156 393790 226208 393796
rect 226064 393780 226116 393786
rect 226064 393722 226116 393728
rect 225972 391740 226024 391746
rect 225972 391682 226024 391688
rect 225708 389146 225920 389174
rect 226352 389174 226380 394318
rect 226628 394176 226656 400044
rect 226444 394148 226656 394176
rect 226444 393718 226472 394148
rect 226720 394074 226748 400044
rect 226536 394046 226748 394074
rect 226432 393712 226484 393718
rect 226432 393654 226484 393660
rect 226352 389146 226472 389174
rect 225604 351416 225656 351422
rect 225604 351358 225656 351364
rect 225512 177608 225564 177614
rect 225512 177550 225564 177556
rect 225420 177540 225472 177546
rect 225420 177482 225472 177488
rect 225328 7948 225380 7954
rect 225328 7890 225380 7896
rect 225144 6180 225196 6186
rect 225144 6122 225196 6128
rect 225708 4146 225736 389146
rect 225696 4140 225748 4146
rect 225696 4082 225748 4088
rect 225052 3936 225104 3942
rect 225052 3878 225104 3884
rect 224224 3732 224276 3738
rect 224224 3674 224276 3680
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 223948 3188 224000 3194
rect 223948 3130 224000 3136
rect 223960 480 223988 3130
rect 225144 2984 225196 2990
rect 225144 2926 225196 2932
rect 225156 480 225184 2926
rect 226352 480 226380 3470
rect 226444 2990 226472 389146
rect 226536 4826 226564 394046
rect 226616 393984 226668 393990
rect 226812 393972 226840 400044
rect 226904 396030 226932 400044
rect 226892 396024 226944 396030
rect 226892 395966 226944 395972
rect 226996 393990 227024 400044
rect 226616 393926 226668 393932
rect 226720 393944 226840 393972
rect 226984 393984 227036 393990
rect 226628 4894 226656 393926
rect 226720 46306 226748 393944
rect 226984 393926 227036 393932
rect 227088 393802 227116 400044
rect 227180 397594 227208 400044
rect 227168 397588 227220 397594
rect 227168 397530 227220 397536
rect 227272 394466 227300 400044
rect 227364 397662 227392 400044
rect 227456 397730 227484 400044
rect 227444 397724 227496 397730
rect 227444 397666 227496 397672
rect 227352 397656 227404 397662
rect 227352 397598 227404 397604
rect 227260 394460 227312 394466
rect 227260 394402 227312 394408
rect 227352 394256 227404 394262
rect 227352 394198 227404 394204
rect 226812 393774 227116 393802
rect 226812 177342 226840 393774
rect 227076 393712 227128 393718
rect 227076 393654 227128 393660
rect 226892 393644 226944 393650
rect 226892 393586 226944 393592
rect 226904 350606 226932 393586
rect 227088 352578 227116 393654
rect 227168 386572 227220 386578
rect 227168 386514 227220 386520
rect 227076 352572 227128 352578
rect 227076 352514 227128 352520
rect 226892 350600 226944 350606
rect 226892 350542 226944 350548
rect 226800 177336 226852 177342
rect 226800 177278 226852 177284
rect 226708 46300 226760 46306
rect 226708 46242 226760 46248
rect 226616 4888 226668 4894
rect 226616 4830 226668 4836
rect 226524 4820 226576 4826
rect 226524 4762 226576 4768
rect 227180 3058 227208 386514
rect 227364 3874 227392 394198
rect 227548 386578 227576 400044
rect 227640 393650 227668 400044
rect 227732 393650 227760 400044
rect 227824 397526 227852 400044
rect 227812 397520 227864 397526
rect 227812 397462 227864 397468
rect 227812 393984 227864 393990
rect 227812 393926 227864 393932
rect 227628 393644 227680 393650
rect 227628 393586 227680 393592
rect 227720 393644 227772 393650
rect 227720 393586 227772 393592
rect 227536 386572 227588 386578
rect 227536 386514 227588 386520
rect 227824 6914 227852 393926
rect 227916 393802 227944 400044
rect 228008 393990 228036 400044
rect 228100 393990 228128 400044
rect 227996 393984 228048 393990
rect 227996 393926 228048 393932
rect 228088 393984 228140 393990
rect 228192 393972 228220 400044
rect 228284 394074 228312 400044
rect 228376 394176 228404 400044
rect 228468 394330 228496 400044
rect 228456 394324 228508 394330
rect 228456 394266 228508 394272
rect 228376 394148 228496 394176
rect 228284 394046 228404 394074
rect 228192 393944 228312 393972
rect 228088 393926 228140 393932
rect 227916 393774 228220 393802
rect 227996 393712 228048 393718
rect 227996 393654 228048 393660
rect 227904 393576 227956 393582
rect 227904 393518 227956 393524
rect 227732 6886 227852 6914
rect 227352 3868 227404 3874
rect 227352 3810 227404 3816
rect 227732 3482 227760 6886
rect 227916 3670 227944 393518
rect 227904 3664 227956 3670
rect 227904 3606 227956 3612
rect 227548 3454 227760 3482
rect 227168 3052 227220 3058
rect 227168 2994 227220 3000
rect 226432 2984 226484 2990
rect 226432 2926 226484 2932
rect 227548 480 227576 3454
rect 228008 3398 228036 393654
rect 228088 393644 228140 393650
rect 228088 393586 228140 393592
rect 227996 3392 228048 3398
rect 227996 3334 228048 3340
rect 228100 3194 228128 393586
rect 228192 3534 228220 393774
rect 228284 3738 228312 393944
rect 228376 393718 228404 394046
rect 228364 393712 228416 393718
rect 228364 393654 228416 393660
rect 228468 393582 228496 394148
rect 228560 394058 228588 400044
rect 228548 394052 228600 394058
rect 228548 393994 228600 394000
rect 228456 393576 228508 393582
rect 228456 393518 228508 393524
rect 228652 389174 228680 400044
rect 228744 397497 228772 400044
rect 228836 397769 228864 400044
rect 228822 397760 228878 397769
rect 228822 397695 228878 397704
rect 228928 397497 228956 400044
rect 229020 397633 229048 400044
rect 229006 397624 229062 397633
rect 229006 397559 229062 397568
rect 228730 397488 228786 397497
rect 228730 397423 228786 397432
rect 228914 397488 228970 397497
rect 228914 397423 228970 397432
rect 228732 394324 228784 394330
rect 228732 394266 228784 394272
rect 228744 391882 228772 394266
rect 228824 393984 228876 393990
rect 228824 393926 228876 393932
rect 228732 391876 228784 391882
rect 228732 391818 228784 391824
rect 228376 389146 228680 389174
rect 228376 352578 228404 389146
rect 228364 352572 228416 352578
rect 228364 352514 228416 352520
rect 228836 6914 228864 393926
rect 229112 392086 229140 400044
rect 229204 392222 229232 400044
rect 229296 393990 229324 400044
rect 229284 393984 229336 393990
rect 229284 393926 229336 393932
rect 229388 393922 229416 400044
rect 229376 393916 229428 393922
rect 229376 393858 229428 393864
rect 229284 393848 229336 393854
rect 229284 393790 229336 393796
rect 229192 392216 229244 392222
rect 229192 392158 229244 392164
rect 229100 392080 229152 392086
rect 229296 392034 229324 393790
rect 229480 392306 229508 400044
rect 229572 393854 229600 400044
rect 229560 393848 229612 393854
rect 229560 393790 229612 393796
rect 229664 392306 229692 400044
rect 229756 398342 229784 400044
rect 229744 398336 229796 398342
rect 229744 398278 229796 398284
rect 229100 392022 229152 392028
rect 228744 6886 228864 6914
rect 229204 392006 229324 392034
rect 229388 392278 229508 392306
rect 229572 392278 229692 392306
rect 228272 3732 228324 3738
rect 228272 3674 228324 3680
rect 228180 3528 228232 3534
rect 228180 3470 228232 3476
rect 228088 3188 228140 3194
rect 228088 3130 228140 3136
rect 228744 480 228772 6886
rect 229204 3874 229232 392006
rect 229284 391944 229336 391950
rect 229284 391886 229336 391892
rect 229192 3868 229244 3874
rect 229192 3810 229244 3816
rect 229296 3602 229324 391886
rect 229284 3596 229336 3602
rect 229284 3538 229336 3544
rect 229388 3466 229416 392278
rect 229468 392216 229520 392222
rect 229468 392158 229520 392164
rect 229480 3942 229508 392158
rect 229572 4894 229600 392278
rect 229848 392170 229876 400044
rect 229664 392142 229876 392170
rect 229560 4888 229612 4894
rect 229560 4830 229612 4836
rect 229664 4826 229692 392142
rect 229744 392080 229796 392086
rect 229744 392022 229796 392028
rect 229756 354074 229784 392022
rect 229940 389174 229968 400044
rect 230032 391950 230060 400044
rect 230124 397497 230152 400044
rect 230216 397905 230244 400044
rect 230202 397896 230258 397905
rect 230202 397831 230258 397840
rect 230308 397769 230336 400044
rect 230294 397760 230350 397769
rect 230294 397695 230350 397704
rect 230400 397633 230428 400044
rect 230386 397624 230442 397633
rect 230386 397559 230442 397568
rect 230110 397488 230166 397497
rect 230110 397423 230166 397432
rect 230492 394074 230520 400044
rect 230584 398274 230612 400044
rect 230572 398268 230624 398274
rect 230572 398210 230624 398216
rect 230400 394046 230520 394074
rect 230112 393984 230164 393990
rect 230112 393926 230164 393932
rect 230020 391944 230072 391950
rect 230020 391886 230072 391892
rect 229848 389146 229968 389174
rect 229744 354068 229796 354074
rect 229744 354010 229796 354016
rect 229848 354006 229876 389146
rect 229836 354000 229888 354006
rect 229836 353942 229888 353948
rect 229652 4820 229704 4826
rect 229652 4762 229704 4768
rect 229468 3936 229520 3942
rect 229468 3878 229520 3884
rect 229836 3732 229888 3738
rect 229836 3674 229888 3680
rect 229376 3460 229428 3466
rect 229376 3402 229428 3408
rect 229848 480 229876 3674
rect 230124 3534 230152 393926
rect 230400 393582 230428 394046
rect 230676 393972 230704 400044
rect 230768 394074 230796 400044
rect 230860 395894 230888 400044
rect 230848 395888 230900 395894
rect 230848 395830 230900 395836
rect 230768 394046 230888 394074
rect 230492 393944 230704 393972
rect 230756 393984 230808 393990
rect 230388 393576 230440 393582
rect 230388 393518 230440 393524
rect 230492 4962 230520 393944
rect 230756 393926 230808 393932
rect 230572 393848 230624 393854
rect 230572 393790 230624 393796
rect 230584 6662 230612 393790
rect 230664 393780 230716 393786
rect 230664 393722 230716 393728
rect 230572 6656 230624 6662
rect 230572 6598 230624 6604
rect 230676 6594 230704 393722
rect 230768 6730 230796 393926
rect 230860 393802 230888 394046
rect 230952 393990 230980 400044
rect 230940 393984 230992 393990
rect 230940 393926 230992 393932
rect 230860 393774 230980 393802
rect 230848 393712 230900 393718
rect 230848 393654 230900 393660
rect 230860 7886 230888 393654
rect 230952 82210 230980 393774
rect 231044 352782 231072 400044
rect 231136 393854 231164 400044
rect 231124 393848 231176 393854
rect 231124 393790 231176 393796
rect 231228 393718 231256 400044
rect 231216 393712 231268 393718
rect 231216 393654 231268 393660
rect 231216 393576 231268 393582
rect 231216 393518 231268 393524
rect 231122 353424 231178 353433
rect 231122 353359 231178 353368
rect 231032 352776 231084 352782
rect 231032 352718 231084 352724
rect 230940 82204 230992 82210
rect 230940 82146 230992 82152
rect 230848 7880 230900 7886
rect 230848 7822 230900 7828
rect 230756 6724 230808 6730
rect 230756 6666 230808 6672
rect 230664 6588 230716 6594
rect 230664 6530 230716 6536
rect 230480 4956 230532 4962
rect 230480 4898 230532 4904
rect 230112 3528 230164 3534
rect 230112 3470 230164 3476
rect 231136 3398 231164 353359
rect 231228 352850 231256 393518
rect 231320 354346 231348 400044
rect 231412 393786 231440 400044
rect 231504 397497 231532 400044
rect 231490 397488 231546 397497
rect 231490 397423 231546 397432
rect 231492 395888 231544 395894
rect 231492 395830 231544 395836
rect 231400 393780 231452 393786
rect 231400 393722 231452 393728
rect 231504 392902 231532 395830
rect 231596 395593 231624 400044
rect 231688 398818 231716 400044
rect 231676 398812 231728 398818
rect 231676 398754 231728 398760
rect 231780 397633 231808 400044
rect 231766 397624 231822 397633
rect 231766 397559 231822 397568
rect 231582 395584 231638 395593
rect 231582 395519 231638 395528
rect 231872 393990 231900 400044
rect 231964 395826 231992 400044
rect 231952 395820 232004 395826
rect 231952 395762 232004 395768
rect 231952 394188 232004 394194
rect 231952 394130 232004 394136
rect 231860 393984 231912 393990
rect 231860 393926 231912 393932
rect 231860 393848 231912 393854
rect 231860 393790 231912 393796
rect 231492 392896 231544 392902
rect 231492 392838 231544 392844
rect 231308 354340 231360 354346
rect 231308 354282 231360 354288
rect 231216 352844 231268 352850
rect 231216 352786 231268 352792
rect 231872 6526 231900 393790
rect 231860 6520 231912 6526
rect 231860 6462 231912 6468
rect 231964 6322 231992 394130
rect 232056 393972 232084 400044
rect 232148 394097 232176 400044
rect 232240 394194 232268 400044
rect 232228 394188 232280 394194
rect 232228 394130 232280 394136
rect 232134 394088 232190 394097
rect 232332 394074 232360 400044
rect 232424 394126 232452 400044
rect 232516 396642 232544 400044
rect 232608 397866 232636 400044
rect 232596 397860 232648 397866
rect 232596 397802 232648 397808
rect 232700 396658 232728 400044
rect 232504 396636 232556 396642
rect 232504 396578 232556 396584
rect 232608 396630 232728 396658
rect 232608 394210 232636 396630
rect 232688 396500 232740 396506
rect 232688 396442 232740 396448
rect 232516 394182 232636 394210
rect 232134 394023 232190 394032
rect 232240 394046 232360 394074
rect 232412 394120 232464 394126
rect 232412 394062 232464 394068
rect 232056 393944 232176 393972
rect 232044 393780 232096 393786
rect 232044 393722 232096 393728
rect 232056 7818 232084 393722
rect 232148 17678 232176 393944
rect 232136 17672 232188 17678
rect 232136 17614 232188 17620
rect 232240 17610 232268 394046
rect 232412 393984 232464 393990
rect 232412 393926 232464 393932
rect 232318 393816 232374 393825
rect 232318 393751 232374 393760
rect 232332 24478 232360 393751
rect 232424 24546 232452 393926
rect 232516 26042 232544 394182
rect 232596 394120 232648 394126
rect 232596 394062 232648 394068
rect 232608 354278 232636 394062
rect 232700 393854 232728 396442
rect 232688 393848 232740 393854
rect 232688 393790 232740 393796
rect 232792 393786 232820 400044
rect 232884 396545 232912 400044
rect 232976 397769 233004 400044
rect 232962 397760 233018 397769
rect 232962 397695 233018 397704
rect 233068 397497 233096 400044
rect 233160 397633 233188 400044
rect 233146 397624 233202 397633
rect 233146 397559 233202 397568
rect 233054 397488 233110 397497
rect 233054 397423 233110 397432
rect 232870 396536 232926 396545
rect 232870 396471 232926 396480
rect 232872 395820 232924 395826
rect 232872 395762 232924 395768
rect 232780 393780 232832 393786
rect 232780 393722 232832 393728
rect 232884 392834 232912 395762
rect 233252 393854 233280 400044
rect 233240 393848 233292 393854
rect 233240 393790 233292 393796
rect 232872 392828 232924 392834
rect 232872 392770 232924 392776
rect 233344 392306 233372 400044
rect 233252 392278 233372 392306
rect 232596 354272 232648 354278
rect 232596 354214 232648 354220
rect 232504 26036 232556 26042
rect 232504 25978 232556 25984
rect 232412 24540 232464 24546
rect 232412 24482 232464 24488
rect 232320 24472 232372 24478
rect 232320 24414 232372 24420
rect 232228 17604 232280 17610
rect 232228 17546 232280 17552
rect 232044 7812 232096 7818
rect 232044 7754 232096 7760
rect 231952 6316 232004 6322
rect 231952 6258 232004 6264
rect 233252 3670 233280 392278
rect 233436 392222 233464 400044
rect 233528 393990 233556 400044
rect 233620 398041 233648 400044
rect 233606 398032 233662 398041
rect 233606 397967 233662 397976
rect 233712 396074 233740 400044
rect 233620 396046 233740 396074
rect 233516 393984 233568 393990
rect 233516 393926 233568 393932
rect 233516 393848 233568 393854
rect 233516 393790 233568 393796
rect 233424 392216 233476 392222
rect 233424 392158 233476 392164
rect 233332 392148 233384 392154
rect 233332 392090 233384 392096
rect 233344 7750 233372 392090
rect 233528 392034 233556 393790
rect 233436 392006 233556 392034
rect 233436 389298 233464 392006
rect 233516 391876 233568 391882
rect 233516 391818 233568 391824
rect 233528 389609 233556 391818
rect 233514 389600 233570 389609
rect 233514 389535 233570 389544
rect 233516 389428 233568 389434
rect 233516 389370 233568 389376
rect 233424 389292 233476 389298
rect 233424 389234 233476 389240
rect 233422 389192 233478 389201
rect 233422 389127 233478 389136
rect 233332 7744 233384 7750
rect 233332 7686 233384 7692
rect 232228 3664 232280 3670
rect 232228 3606 232280 3612
rect 233240 3664 233292 3670
rect 233240 3606 233292 3612
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231124 3392 231176 3398
rect 231124 3334 231176 3340
rect 231044 480 231072 3334
rect 232240 480 232268 3606
rect 233436 480 233464 389127
rect 233528 18970 233556 389370
rect 233620 19038 233648 396046
rect 233804 394330 233832 400044
rect 233792 394324 233844 394330
rect 233792 394266 233844 394272
rect 233792 393984 233844 393990
rect 233792 393926 233844 393932
rect 233700 392216 233752 392222
rect 233700 392158 233752 392164
rect 233712 19106 233740 392158
rect 233804 389314 233832 393926
rect 233896 392154 233924 400044
rect 233884 392148 233936 392154
rect 233884 392090 233936 392096
rect 233988 389434 234016 400044
rect 234080 397497 234108 400044
rect 234172 397633 234200 400044
rect 234158 397624 234214 397633
rect 234158 397559 234214 397568
rect 234066 397488 234122 397497
rect 234066 397423 234122 397432
rect 234264 397186 234292 400044
rect 234252 397180 234304 397186
rect 234252 397122 234304 397128
rect 234356 394466 234384 400044
rect 234448 397769 234476 400044
rect 234434 397760 234490 397769
rect 234434 397695 234490 397704
rect 234540 397497 234568 400044
rect 234526 397488 234582 397497
rect 234526 397423 234582 397432
rect 234344 394460 234396 394466
rect 234344 394402 234396 394408
rect 234068 394324 234120 394330
rect 234068 394266 234120 394272
rect 234080 389842 234108 394266
rect 234632 394194 234660 400044
rect 234724 397594 234752 400044
rect 234712 397588 234764 397594
rect 234712 397530 234764 397536
rect 234712 394324 234764 394330
rect 234712 394266 234764 394272
rect 234620 394188 234672 394194
rect 234620 394130 234672 394136
rect 234620 394052 234672 394058
rect 234620 393994 234672 394000
rect 234160 393916 234212 393922
rect 234160 393858 234212 393864
rect 234068 389836 234120 389842
rect 234068 389778 234120 389784
rect 233976 389428 234028 389434
rect 233976 389370 234028 389376
rect 233804 389286 234016 389314
rect 233792 389224 233844 389230
rect 233792 389166 233844 389172
rect 233884 389224 233936 389230
rect 233884 389166 233936 389172
rect 233804 177750 233832 389166
rect 233792 177744 233844 177750
rect 233792 177686 233844 177692
rect 233700 19100 233752 19106
rect 233700 19042 233752 19048
rect 233608 19032 233660 19038
rect 233608 18974 233660 18980
rect 233516 18964 233568 18970
rect 233516 18906 233568 18912
rect 233896 4010 233924 389166
rect 233988 177682 234016 389286
rect 234172 389230 234200 393858
rect 234160 389224 234212 389230
rect 234160 389166 234212 389172
rect 233976 177676 234028 177682
rect 233976 177618 234028 177624
rect 233884 4004 233936 4010
rect 233884 3946 233936 3952
rect 234632 480 234660 393994
rect 234724 9450 234752 394266
rect 234816 18902 234844 400044
rect 234908 393825 234936 400044
rect 235000 394126 235028 400044
rect 234988 394120 235040 394126
rect 234988 394062 235040 394068
rect 234894 393816 234950 393825
rect 235092 393802 235120 400044
rect 235184 394398 235212 400044
rect 235172 394392 235224 394398
rect 235172 394334 235224 394340
rect 235276 394330 235304 400044
rect 235264 394324 235316 394330
rect 235264 394266 235316 394272
rect 235368 394210 235396 400044
rect 235172 394188 235224 394194
rect 235172 394130 235224 394136
rect 235276 394182 235396 394210
rect 234894 393751 234950 393760
rect 235000 393774 235120 393802
rect 234896 393712 234948 393718
rect 234896 393654 234948 393660
rect 234804 18896 234856 18902
rect 234804 18838 234856 18844
rect 234908 18766 234936 393654
rect 235000 18834 235028 393774
rect 235080 393712 235132 393718
rect 235080 393654 235132 393660
rect 235092 25906 235120 393654
rect 235184 25974 235212 394130
rect 235276 393922 235304 394182
rect 235356 394120 235408 394126
rect 235356 394062 235408 394068
rect 235264 393916 235316 393922
rect 235264 393858 235316 393864
rect 235262 393816 235318 393825
rect 235262 393751 235318 393760
rect 235276 355706 235304 393751
rect 235264 355700 235316 355706
rect 235264 355642 235316 355648
rect 235264 352572 235316 352578
rect 235264 352514 235316 352520
rect 235172 25968 235224 25974
rect 235172 25910 235224 25916
rect 235080 25900 235132 25906
rect 235080 25842 235132 25848
rect 234988 18828 235040 18834
rect 234988 18770 235040 18776
rect 234896 18760 234948 18766
rect 234896 18702 234948 18708
rect 235276 16574 235304 352514
rect 235368 87786 235396 394062
rect 235460 393718 235488 400044
rect 235448 393712 235500 393718
rect 235448 393654 235500 393660
rect 235552 389174 235580 400044
rect 235644 397225 235672 400044
rect 235736 397633 235764 400044
rect 235722 397624 235778 397633
rect 235722 397559 235778 397568
rect 235828 397497 235856 400044
rect 235814 397488 235870 397497
rect 235814 397423 235870 397432
rect 235630 397216 235686 397225
rect 235630 397151 235686 397160
rect 235920 397089 235948 400044
rect 235906 397080 235962 397089
rect 235906 397015 235962 397024
rect 236012 394670 236040 400044
rect 236104 398546 236132 400044
rect 236092 398540 236144 398546
rect 236092 398482 236144 398488
rect 236000 394664 236052 394670
rect 236000 394606 236052 394612
rect 236000 394052 236052 394058
rect 236000 393994 236052 394000
rect 235460 389146 235580 389174
rect 235460 355638 235488 389146
rect 235448 355632 235500 355638
rect 235448 355574 235500 355580
rect 235356 87780 235408 87786
rect 235356 87722 235408 87728
rect 235276 16546 235856 16574
rect 234712 9444 234764 9450
rect 234712 9386 234764 9392
rect 235828 480 235856 16546
rect 236012 9314 236040 393994
rect 236092 393984 236144 393990
rect 236092 393926 236144 393932
rect 236104 9382 236132 393926
rect 236196 18698 236224 400044
rect 236288 393972 236316 400044
rect 236380 398682 236408 400044
rect 236368 398676 236420 398682
rect 236368 398618 236420 398624
rect 236288 393944 236408 393972
rect 236276 393508 236328 393514
rect 236276 393450 236328 393456
rect 236184 18692 236236 18698
rect 236184 18634 236236 18640
rect 236288 18630 236316 393450
rect 236380 391338 236408 393944
rect 236472 393514 236500 400044
rect 236460 393508 236512 393514
rect 236460 393450 236512 393456
rect 236564 391354 236592 400044
rect 236656 393990 236684 400044
rect 236748 396846 236776 400044
rect 236736 396840 236788 396846
rect 236736 396782 236788 396788
rect 236840 394602 236868 400044
rect 236828 394596 236880 394602
rect 236828 394538 236880 394544
rect 236932 394058 236960 400044
rect 236920 394052 236972 394058
rect 236920 393994 236972 394000
rect 236644 393984 236696 393990
rect 236644 393926 236696 393932
rect 236368 391332 236420 391338
rect 236368 391274 236420 391280
rect 236472 391326 236592 391354
rect 236472 391218 236500 391326
rect 236380 391190 236500 391218
rect 236380 23186 236408 391190
rect 236460 391128 236512 391134
rect 236460 391070 236512 391076
rect 236472 25838 236500 391070
rect 237024 389174 237052 400044
rect 237116 397497 237144 400044
rect 237208 397769 237236 400044
rect 237194 397760 237250 397769
rect 237194 397695 237250 397704
rect 237300 397633 237328 400044
rect 237286 397624 237342 397633
rect 237286 397559 237342 397568
rect 237102 397488 237158 397497
rect 237102 397423 237158 397432
rect 237392 397338 237420 400044
rect 237484 397458 237512 400044
rect 237472 397452 237524 397458
rect 237472 397394 237524 397400
rect 237392 397310 237512 397338
rect 237380 397180 237432 397186
rect 237380 397122 237432 397128
rect 236564 389146 237052 389174
rect 236564 351286 236592 389146
rect 236642 353560 236698 353569
rect 236642 353495 236698 353504
rect 236552 351280 236604 351286
rect 236552 351222 236604 351228
rect 236460 25832 236512 25838
rect 236460 25774 236512 25780
rect 236368 23180 236420 23186
rect 236368 23122 236420 23128
rect 236276 18624 236328 18630
rect 236276 18566 236328 18572
rect 236092 9376 236144 9382
rect 236092 9318 236144 9324
rect 236000 9308 236052 9314
rect 236000 9250 236052 9256
rect 236656 3670 236684 353495
rect 237392 5166 237420 397122
rect 237484 394534 237512 397310
rect 237472 394528 237524 394534
rect 237472 394470 237524 394476
rect 237472 393984 237524 393990
rect 237472 393926 237524 393932
rect 237484 9178 237512 393926
rect 237576 392222 237604 400044
rect 237668 397050 237696 400044
rect 237656 397044 237708 397050
rect 237656 396986 237708 396992
rect 237760 392306 237788 400044
rect 237668 392278 237788 392306
rect 237564 392216 237616 392222
rect 237564 392158 237616 392164
rect 237564 392080 237616 392086
rect 237564 392022 237616 392028
rect 237472 9172 237524 9178
rect 237472 9114 237524 9120
rect 237576 9110 237604 392022
rect 237668 9246 237696 392278
rect 237748 392216 237800 392222
rect 237748 392158 237800 392164
rect 237760 20262 237788 392158
rect 237748 20256 237800 20262
rect 237748 20198 237800 20204
rect 237852 20194 237880 400044
rect 237944 397186 237972 400044
rect 237932 397180 237984 397186
rect 237932 397122 237984 397128
rect 237932 397044 237984 397050
rect 237932 396986 237984 396992
rect 237944 356726 237972 396986
rect 238036 393990 238064 400044
rect 238024 393984 238076 393990
rect 238024 393926 238076 393932
rect 238128 389174 238156 400044
rect 238220 397526 238248 400044
rect 238208 397520 238260 397526
rect 238208 397462 238260 397468
rect 238312 392086 238340 400044
rect 238404 397633 238432 400044
rect 238496 397769 238524 400044
rect 238482 397760 238538 397769
rect 238482 397695 238538 397704
rect 238390 397624 238446 397633
rect 238390 397559 238446 397568
rect 238588 397497 238616 400044
rect 238574 397488 238630 397497
rect 238392 397452 238444 397458
rect 238574 397423 238630 397432
rect 238392 397394 238444 397400
rect 238404 392766 238432 397394
rect 238680 396953 238708 400044
rect 238772 397866 238800 400044
rect 238760 397860 238812 397866
rect 238760 397802 238812 397808
rect 238666 396944 238722 396953
rect 238666 396879 238722 396888
rect 238760 393984 238812 393990
rect 238864 393972 238892 400044
rect 238956 394074 238984 400044
rect 239048 394194 239076 400044
rect 239036 394188 239088 394194
rect 239036 394130 239088 394136
rect 238956 394046 239076 394074
rect 238864 393944 238984 393972
rect 238760 393926 238812 393932
rect 238392 392760 238444 392766
rect 238392 392702 238444 392708
rect 238300 392080 238352 392086
rect 238300 392022 238352 392028
rect 238036 389146 238156 389174
rect 237932 356720 237984 356726
rect 237932 356662 237984 356668
rect 238036 354210 238064 389146
rect 238024 354204 238076 354210
rect 238024 354146 238076 354152
rect 237930 353968 237986 353977
rect 237930 353903 237986 353912
rect 237840 20188 237892 20194
rect 237840 20130 237892 20136
rect 237656 9240 237708 9246
rect 237656 9182 237708 9188
rect 237564 9104 237616 9110
rect 237564 9046 237616 9052
rect 237380 5160 237432 5166
rect 237380 5102 237432 5108
rect 236644 3664 236696 3670
rect 236644 3606 236696 3612
rect 237012 3392 237064 3398
rect 237012 3334 237064 3340
rect 237024 480 237052 3334
rect 220004 354 220032 462
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237944 354 237972 353903
rect 238772 10538 238800 393926
rect 238852 393848 238904 393854
rect 238852 393790 238904 393796
rect 238864 10606 238892 393790
rect 238956 10674 238984 393944
rect 239048 393700 239076 394046
rect 239140 393854 239168 400044
rect 239232 393972 239260 400044
rect 239324 397798 239352 400044
rect 239312 397792 239364 397798
rect 239312 397734 239364 397740
rect 239416 393990 239444 400044
rect 239404 393984 239456 393990
rect 239232 393944 239352 393972
rect 239128 393848 239180 393854
rect 239128 393790 239180 393796
rect 239048 393672 239260 393700
rect 239128 393576 239180 393582
rect 239128 393518 239180 393524
rect 239036 393508 239088 393514
rect 239036 393450 239088 393456
rect 239048 20126 239076 393450
rect 239140 25770 239168 393518
rect 239232 355502 239260 393672
rect 239220 355496 239272 355502
rect 239220 355438 239272 355444
rect 239324 355434 239352 393944
rect 239404 393926 239456 393932
rect 239508 393514 239536 400044
rect 239600 393582 239628 400044
rect 239692 397769 239720 400044
rect 239678 397760 239734 397769
rect 239678 397695 239734 397704
rect 239680 397656 239732 397662
rect 239784 397633 239812 400044
rect 239876 397662 239904 400044
rect 239864 397656 239916 397662
rect 239680 397598 239732 397604
rect 239770 397624 239826 397633
rect 239588 393576 239640 393582
rect 239588 393518 239640 393524
rect 239496 393508 239548 393514
rect 239496 393450 239548 393456
rect 239692 389174 239720 397598
rect 239864 397598 239916 397604
rect 239770 397559 239826 397568
rect 239968 397497 239996 400044
rect 240060 397905 240088 400044
rect 240046 397896 240102 397905
rect 240046 397831 240102 397840
rect 240048 397588 240100 397594
rect 240048 397530 240100 397536
rect 239954 397488 240010 397497
rect 239954 397423 240010 397432
rect 240060 391542 240088 397530
rect 240152 394330 240180 400044
rect 240244 399022 240272 400044
rect 240232 399016 240284 399022
rect 240232 398958 240284 398964
rect 240336 395146 240364 400044
rect 240428 397730 240456 400044
rect 240416 397724 240468 397730
rect 240416 397666 240468 397672
rect 240324 395140 240376 395146
rect 240324 395082 240376 395088
rect 240140 394324 240192 394330
rect 240140 394266 240192 394272
rect 240520 394074 240548 400044
rect 240152 394046 240548 394074
rect 240048 391536 240100 391542
rect 240048 391478 240100 391484
rect 239416 389146 239720 389174
rect 239312 355428 239364 355434
rect 239312 355370 239364 355376
rect 239416 84930 239444 389146
rect 239404 84924 239456 84930
rect 239404 84866 239456 84872
rect 239128 25764 239180 25770
rect 239128 25706 239180 25712
rect 239036 20120 239088 20126
rect 239036 20062 239088 20068
rect 238944 10668 238996 10674
rect 238944 10610 238996 10616
rect 238852 10600 238904 10606
rect 238852 10542 238904 10548
rect 238760 10532 238812 10538
rect 238760 10474 238812 10480
rect 240152 10470 240180 394046
rect 240416 393984 240468 393990
rect 240612 393972 240640 400044
rect 240416 393926 240468 393932
rect 240520 393944 240640 393972
rect 240232 393916 240284 393922
rect 240232 393858 240284 393864
rect 240140 10464 240192 10470
rect 240140 10406 240192 10412
rect 240244 10402 240272 393858
rect 240324 393848 240376 393854
rect 240324 393790 240376 393796
rect 240336 12102 240364 393790
rect 240428 19990 240456 393926
rect 240520 20058 240548 393944
rect 240704 393904 240732 400044
rect 240796 393922 240824 400044
rect 240888 393990 240916 400044
rect 240980 397594 241008 400044
rect 240968 397588 241020 397594
rect 240968 397530 241020 397536
rect 240968 395140 241020 395146
rect 240968 395082 241020 395088
rect 240876 393984 240928 393990
rect 240876 393926 240928 393932
rect 240612 393876 240732 393904
rect 240784 393916 240836 393922
rect 240612 177546 240640 393876
rect 240784 393858 240836 393864
rect 240980 391474 241008 395082
rect 241072 393854 241100 400044
rect 241164 396778 241192 400044
rect 241152 396772 241204 396778
rect 241152 396714 241204 396720
rect 241152 394324 241204 394330
rect 241152 394266 241204 394272
rect 241060 393848 241112 393854
rect 241060 393790 241112 393796
rect 240968 391468 241020 391474
rect 240968 391410 241020 391416
rect 241164 391218 241192 394266
rect 240704 391190 241192 391218
rect 240704 177614 240732 391190
rect 241256 389174 241284 400044
rect 241348 397497 241376 400044
rect 241440 397633 241468 400044
rect 241532 398954 241560 400044
rect 241520 398948 241572 398954
rect 241520 398890 241572 398896
rect 241426 397624 241482 397633
rect 241426 397559 241482 397568
rect 241334 397488 241390 397497
rect 241334 397423 241390 397432
rect 241520 394324 241572 394330
rect 241520 394266 241572 394272
rect 240796 389146 241284 389174
rect 240796 354142 240824 389146
rect 240784 354136 240836 354142
rect 240784 354078 240836 354084
rect 240692 177608 240744 177614
rect 240692 177550 240744 177556
rect 240600 177540 240652 177546
rect 240600 177482 240652 177488
rect 240508 20052 240560 20058
rect 240508 19994 240560 20000
rect 240416 19984 240468 19990
rect 240416 19926 240468 19932
rect 240324 12096 240376 12102
rect 240324 12038 240376 12044
rect 240232 10396 240284 10402
rect 240232 10338 240284 10344
rect 241532 6458 241560 394266
rect 241624 394074 241652 400044
rect 241716 394194 241744 400044
rect 241808 394330 241836 400044
rect 241796 394324 241848 394330
rect 241796 394266 241848 394272
rect 241704 394188 241756 394194
rect 241704 394130 241756 394136
rect 241624 394046 241744 394074
rect 241612 393848 241664 393854
rect 241612 393790 241664 393796
rect 241520 6452 241572 6458
rect 241520 6394 241572 6400
rect 241624 6390 241652 393790
rect 241716 12034 241744 394046
rect 241796 393984 241848 393990
rect 241796 393926 241848 393932
rect 241704 12028 241756 12034
rect 241704 11970 241756 11976
rect 241808 11898 241836 393926
rect 241900 11966 241928 400044
rect 241992 394058 242020 400044
rect 242084 398138 242112 400044
rect 242072 398132 242124 398138
rect 242072 398074 242124 398080
rect 242176 396642 242204 400044
rect 242164 396636 242216 396642
rect 242164 396578 242216 396584
rect 242268 394346 242296 400044
rect 242360 396522 242388 400044
rect 242452 397769 242480 400044
rect 242438 397760 242494 397769
rect 242438 397695 242494 397704
rect 242544 397633 242572 400044
rect 242636 398886 242664 400044
rect 242624 398880 242676 398886
rect 242624 398822 242676 398828
rect 242622 398712 242678 398721
rect 242622 398647 242678 398656
rect 242530 397624 242586 397633
rect 242530 397559 242586 397568
rect 242532 397520 242584 397526
rect 242532 397462 242584 397468
rect 242360 396494 242480 396522
rect 242348 396432 242400 396438
rect 242348 396374 242400 396380
rect 242084 394318 242296 394346
rect 241980 394052 242032 394058
rect 241980 393994 242032 394000
rect 242084 389174 242112 394318
rect 242164 394188 242216 394194
rect 242164 394130 242216 394136
rect 241992 389146 242112 389174
rect 241992 21894 242020 389146
rect 242072 354068 242124 354074
rect 242072 354010 242124 354016
rect 241980 21888 242032 21894
rect 241980 21830 242032 21836
rect 241888 11960 241940 11966
rect 241888 11902 241940 11908
rect 241796 11892 241848 11898
rect 241796 11834 241848 11840
rect 241612 6384 241664 6390
rect 241612 6326 241664 6332
rect 239404 4956 239456 4962
rect 239404 4898 239456 4904
rect 239416 3874 239444 4898
rect 239220 3868 239272 3874
rect 239220 3810 239272 3816
rect 239404 3868 239456 3874
rect 239404 3810 239456 3816
rect 239232 3398 239260 3810
rect 239310 3496 239366 3505
rect 239310 3431 239366 3440
rect 239220 3392 239272 3398
rect 239220 3334 239272 3340
rect 239324 480 239352 3431
rect 240506 3360 240562 3369
rect 240506 3295 240562 3304
rect 240520 480 240548 3295
rect 238086 354 238198 480
rect 237944 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 354010
rect 242176 83502 242204 394130
rect 242256 394052 242308 394058
rect 242256 393994 242308 394000
rect 242268 87718 242296 393994
rect 242360 393990 242388 396374
rect 242348 393984 242400 393990
rect 242348 393926 242400 393932
rect 242452 393854 242480 396494
rect 242440 393848 242492 393854
rect 242440 393790 242492 393796
rect 242544 389174 242572 397462
rect 242636 396817 242664 398647
rect 242728 397497 242756 400044
rect 242820 398993 242848 400044
rect 242806 398984 242862 398993
rect 242806 398919 242862 398928
rect 242808 398880 242860 398886
rect 242808 398822 242860 398828
rect 242820 398614 242848 398822
rect 242808 398608 242860 398614
rect 242808 398550 242860 398556
rect 242808 397860 242860 397866
rect 242808 397802 242860 397808
rect 242714 397488 242770 397497
rect 242714 397423 242770 397432
rect 242820 397168 242848 397802
rect 242728 397140 242848 397168
rect 242622 396808 242678 396817
rect 242622 396743 242678 396752
rect 242728 394126 242756 397140
rect 242912 394330 242940 400044
rect 243004 395146 243032 400044
rect 242992 395140 243044 395146
rect 242992 395082 243044 395088
rect 243096 394516 243124 400044
rect 243188 397526 243216 400044
rect 243176 397520 243228 397526
rect 243176 397462 243228 397468
rect 243004 394488 243124 394516
rect 243004 394346 243032 394488
rect 242900 394324 242952 394330
rect 243004 394318 243124 394346
rect 242900 394266 242952 394272
rect 242808 394256 242860 394262
rect 242808 394198 242860 394204
rect 242716 394120 242768 394126
rect 242716 394062 242768 394068
rect 242820 393972 242848 394198
rect 242992 393984 243044 393990
rect 242820 393944 242940 393972
rect 242452 389146 242572 389174
rect 242452 355570 242480 389146
rect 242440 355564 242492 355570
rect 242440 355506 242492 355512
rect 242256 87712 242308 87718
rect 242256 87654 242308 87660
rect 242164 83496 242216 83502
rect 242164 83438 242216 83444
rect 242912 11762 242940 393944
rect 242992 393926 243044 393932
rect 243004 11830 243032 393926
rect 243096 393854 243124 394318
rect 243176 394324 243228 394330
rect 243176 394266 243228 394272
rect 243084 393848 243136 393854
rect 243084 393790 243136 393796
rect 243084 393712 243136 393718
rect 243084 393654 243136 393660
rect 243096 13530 243124 393654
rect 243188 16318 243216 394266
rect 243280 393990 243308 400044
rect 243268 393984 243320 393990
rect 243268 393926 243320 393932
rect 243268 393780 243320 393786
rect 243268 393722 243320 393728
rect 243280 21690 243308 393722
rect 243372 21758 243400 400044
rect 243464 393972 243492 400044
rect 243556 394262 243584 400044
rect 243544 394256 243596 394262
rect 243544 394198 243596 394204
rect 243464 393944 243584 393972
rect 243452 393848 243504 393854
rect 243452 393790 243504 393796
rect 243464 21826 243492 393790
rect 243556 25702 243584 393944
rect 243648 393786 243676 400044
rect 243740 398274 243768 400044
rect 243728 398268 243780 398274
rect 243728 398210 243780 398216
rect 243728 395140 243780 395146
rect 243728 395082 243780 395088
rect 243636 393780 243688 393786
rect 243636 393722 243688 393728
rect 243740 391406 243768 395082
rect 243832 393718 243860 400044
rect 243924 397905 243952 400044
rect 243910 397896 243966 397905
rect 243910 397831 243966 397840
rect 244016 397769 244044 400044
rect 244002 397760 244058 397769
rect 244002 397695 244058 397704
rect 243912 397656 243964 397662
rect 243912 397598 243964 397604
rect 243924 393990 243952 397598
rect 244108 397497 244136 400044
rect 244200 397633 244228 400044
rect 244292 398750 244320 400044
rect 244280 398744 244332 398750
rect 244280 398686 244332 398692
rect 244186 397624 244242 397633
rect 244186 397559 244242 397568
rect 244094 397488 244150 397497
rect 244094 397423 244150 397432
rect 244384 397202 244412 400044
rect 244200 397174 244412 397202
rect 244200 396166 244228 397174
rect 244188 396160 244240 396166
rect 244188 396102 244240 396108
rect 244188 394664 244240 394670
rect 244188 394606 244240 394612
rect 244096 394596 244148 394602
rect 244096 394538 244148 394544
rect 244004 394528 244056 394534
rect 244004 394470 244056 394476
rect 244016 394194 244044 394470
rect 244108 394262 244136 394538
rect 244200 394330 244228 394606
rect 244372 394596 244424 394602
rect 244372 394538 244424 394544
rect 244280 394528 244332 394534
rect 244280 394470 244332 394476
rect 244188 394324 244240 394330
rect 244188 394266 244240 394272
rect 244096 394256 244148 394262
rect 244096 394198 244148 394204
rect 244004 394188 244056 394194
rect 244004 394130 244056 394136
rect 243912 393984 243964 393990
rect 243912 393926 243964 393932
rect 243820 393712 243872 393718
rect 243820 393654 243872 393660
rect 243728 391400 243780 391406
rect 243728 391342 243780 391348
rect 243544 25696 243596 25702
rect 243544 25638 243596 25644
rect 243452 21820 243504 21826
rect 243452 21762 243504 21768
rect 243360 21752 243412 21758
rect 243360 21694 243412 21700
rect 243268 21684 243320 21690
rect 243268 21626 243320 21632
rect 243176 16312 243228 16318
rect 243176 16254 243228 16260
rect 243084 13524 243136 13530
rect 243084 13466 243136 13472
rect 244292 13462 244320 394470
rect 244384 393802 244412 394538
rect 244476 393972 244504 400044
rect 244568 394670 244596 400044
rect 244556 394664 244608 394670
rect 244556 394606 244608 394612
rect 244660 394534 244688 400044
rect 244648 394528 244700 394534
rect 244648 394470 244700 394476
rect 244476 393944 244596 393972
rect 244384 393774 244504 393802
rect 244372 393712 244424 393718
rect 244372 393654 244424 393660
rect 244280 13456 244332 13462
rect 244280 13398 244332 13404
rect 244384 13326 244412 393654
rect 244476 13394 244504 393774
rect 244568 21622 244596 393944
rect 244752 393768 244780 400044
rect 244844 397662 244872 400044
rect 244832 397656 244884 397662
rect 244832 397598 244884 397604
rect 244832 394664 244884 394670
rect 244832 394606 244884 394612
rect 244844 394482 244872 394606
rect 244936 394602 244964 400044
rect 244924 394596 244976 394602
rect 244924 394538 244976 394544
rect 244844 394454 244964 394482
rect 244660 393740 244780 393768
rect 244556 21616 244608 21622
rect 244556 21558 244608 21564
rect 244660 21554 244688 393740
rect 244936 393530 244964 394454
rect 244752 393502 244964 393530
rect 244752 25634 244780 393502
rect 245028 392698 245056 400044
rect 245016 392692 245068 392698
rect 245016 392634 245068 392640
rect 245120 392578 245148 400044
rect 245212 393718 245240 400044
rect 245200 393712 245252 393718
rect 245200 393654 245252 393660
rect 244844 392550 245148 392578
rect 244740 25628 244792 25634
rect 244740 25570 244792 25576
rect 244844 25566 244872 392550
rect 245304 389174 245332 400044
rect 245396 399129 245424 400044
rect 245382 399120 245438 399129
rect 245382 399055 245438 399064
rect 245488 397497 245516 400044
rect 245580 397633 245608 400044
rect 245672 397866 245700 400044
rect 245764 398886 245792 400044
rect 245752 398880 245804 398886
rect 245752 398822 245804 398828
rect 245660 397860 245712 397866
rect 245660 397802 245712 397808
rect 245566 397624 245622 397633
rect 245566 397559 245622 397568
rect 245474 397488 245530 397497
rect 245474 397423 245530 397432
rect 245384 396160 245436 396166
rect 245384 396102 245436 396108
rect 245396 391338 245424 396102
rect 245856 396074 245884 400044
rect 245948 397322 245976 400044
rect 245936 397316 245988 397322
rect 245936 397258 245988 397264
rect 245856 396046 245976 396074
rect 245752 394528 245804 394534
rect 245752 394470 245804 394476
rect 245660 393916 245712 393922
rect 245660 393858 245712 393864
rect 245384 391332 245436 391338
rect 245384 391274 245436 391280
rect 244936 389146 245332 389174
rect 244936 87650 244964 389146
rect 244924 87644 244976 87650
rect 244924 87586 244976 87592
rect 244832 25560 244884 25566
rect 244832 25502 244884 25508
rect 244648 21548 244700 21554
rect 244648 21490 244700 21496
rect 244464 13388 244516 13394
rect 244464 13330 244516 13336
rect 244372 13320 244424 13326
rect 244372 13262 244424 13268
rect 245672 13190 245700 393858
rect 245764 13258 245792 394470
rect 245948 394346 245976 396046
rect 246040 394534 246068 400044
rect 246028 394528 246080 394534
rect 246028 394470 246080 394476
rect 245948 394318 246068 394346
rect 245844 393848 245896 393854
rect 245844 393790 245896 393796
rect 245752 13252 245804 13258
rect 245752 13194 245804 13200
rect 245660 13184 245712 13190
rect 245660 13126 245712 13132
rect 245856 13122 245884 393790
rect 245936 393780 245988 393786
rect 245936 393722 245988 393728
rect 245948 21418 245976 393722
rect 246040 21486 246068 394318
rect 246132 393786 246160 400044
rect 246224 397934 246252 400044
rect 246212 397928 246264 397934
rect 246212 397870 246264 397876
rect 246212 397724 246264 397730
rect 246212 397666 246264 397672
rect 246120 393780 246172 393786
rect 246120 393722 246172 393728
rect 246120 393644 246172 393650
rect 246120 393586 246172 393592
rect 246132 23118 246160 393586
rect 246224 389174 246252 397666
rect 246316 393922 246344 400044
rect 246304 393916 246356 393922
rect 246304 393858 246356 393864
rect 246408 393650 246436 400044
rect 246500 397497 246528 400044
rect 246486 397488 246542 397497
rect 246486 397423 246542 397432
rect 246592 393854 246620 400044
rect 246684 397633 246712 400044
rect 246776 398478 246804 400044
rect 246764 398472 246816 398478
rect 246764 398414 246816 398420
rect 246764 397792 246816 397798
rect 246764 397734 246816 397740
rect 246670 397624 246726 397633
rect 246670 397559 246726 397568
rect 246776 395758 246804 397734
rect 246868 397497 246896 400044
rect 246960 397769 246988 400044
rect 246946 397760 247002 397769
rect 246946 397695 247002 397704
rect 246948 397588 247000 397594
rect 246948 397530 247000 397536
rect 246854 397488 246910 397497
rect 246854 397423 246910 397432
rect 246764 395752 246816 395758
rect 246764 395694 246816 395700
rect 246580 393848 246632 393854
rect 246580 393790 246632 393796
rect 246396 393644 246448 393650
rect 246396 393586 246448 393592
rect 246960 389174 246988 397530
rect 247052 394670 247080 400044
rect 247040 394664 247092 394670
rect 247040 394606 247092 394612
rect 246224 389146 246344 389174
rect 246316 228410 246344 389146
rect 246684 389146 246988 389174
rect 246684 355366 246712 389146
rect 246672 355360 246724 355366
rect 246672 355302 246724 355308
rect 246304 228404 246356 228410
rect 246304 228346 246356 228352
rect 246120 23112 246172 23118
rect 246120 23054 246172 23060
rect 246028 21480 246080 21486
rect 246028 21422 246080 21428
rect 245936 21412 245988 21418
rect 245936 21354 245988 21360
rect 247144 14822 247172 400044
rect 247236 393922 247264 400044
rect 247328 398449 247356 400044
rect 247314 398440 247370 398449
rect 247314 398375 247370 398384
rect 247224 393916 247276 393922
rect 247224 393858 247276 393864
rect 247420 393802 247448 400044
rect 247236 393774 247448 393802
rect 247132 14816 247184 14822
rect 247132 14758 247184 14764
rect 247236 14754 247264 393774
rect 247408 393712 247460 393718
rect 247408 393654 247460 393660
rect 247316 390448 247368 390454
rect 247316 390390 247368 390396
rect 247224 14748 247276 14754
rect 247224 14690 247276 14696
rect 247328 14686 247356 390390
rect 247420 23050 247448 393654
rect 247512 82142 247540 400044
rect 247604 390386 247632 400044
rect 247696 395690 247724 400044
rect 247684 395684 247736 395690
rect 247684 395626 247736 395632
rect 247788 390454 247816 400044
rect 247776 390448 247828 390454
rect 247776 390390 247828 390396
rect 247592 390380 247644 390386
rect 247592 390322 247644 390328
rect 247880 390266 247908 400044
rect 247604 390238 247908 390266
rect 247604 86358 247632 390238
rect 247776 390176 247828 390182
rect 247776 390118 247828 390124
rect 247788 386414 247816 390118
rect 247972 389174 248000 400044
rect 248064 397497 248092 400044
rect 248156 397769 248184 400044
rect 248142 397760 248198 397769
rect 248142 397695 248198 397704
rect 248248 397497 248276 400044
rect 248340 397633 248368 400044
rect 248326 397624 248382 397633
rect 248326 397559 248382 397568
rect 248050 397488 248106 397497
rect 248050 397423 248106 397432
rect 248234 397488 248290 397497
rect 248234 397423 248290 397432
rect 248052 395684 248104 395690
rect 248052 395626 248104 395632
rect 248064 392630 248092 395626
rect 248432 393922 248460 400044
rect 248524 398177 248552 400044
rect 248510 398168 248566 398177
rect 248510 398103 248566 398112
rect 248616 393972 248644 400044
rect 248708 395078 248736 400044
rect 248800 398585 248828 400044
rect 248786 398576 248842 398585
rect 248786 398511 248842 398520
rect 248696 395072 248748 395078
rect 248696 395014 248748 395020
rect 248892 394074 248920 400044
rect 248524 393944 248644 393972
rect 248708 394046 248920 394074
rect 248420 393916 248472 393922
rect 248420 393858 248472 393864
rect 248420 393780 248472 393786
rect 248420 393722 248472 393728
rect 248052 392624 248104 392630
rect 248052 392566 248104 392572
rect 247972 389146 248092 389174
rect 247696 386386 247816 386414
rect 247696 177478 247724 386386
rect 247684 177472 247736 177478
rect 247684 177414 247736 177420
rect 247592 86352 247644 86358
rect 247592 86294 247644 86300
rect 247500 82136 247552 82142
rect 247500 82078 247552 82084
rect 247408 23044 247460 23050
rect 247408 22986 247460 22992
rect 247316 14680 247368 14686
rect 247316 14622 247368 14628
rect 245844 13116 245896 13122
rect 245844 13058 245896 13064
rect 242992 11824 243044 11830
rect 242992 11766 243044 11772
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 245200 4004 245252 4010
rect 245200 3946 245252 3952
rect 242900 3936 242952 3942
rect 242900 3878 242952 3884
rect 242912 480 242940 3878
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 244108 480 244136 3470
rect 245212 480 245240 3946
rect 248064 3534 248092 389146
rect 248432 5098 248460 393722
rect 248524 14618 248552 393944
rect 248708 393802 248736 394046
rect 248984 393972 249012 400044
rect 248892 393944 249012 393972
rect 248788 393916 248840 393922
rect 248788 393858 248840 393864
rect 248616 393774 248736 393802
rect 248512 14612 248564 14618
rect 248512 14554 248564 14560
rect 248616 14550 248644 393774
rect 248696 393712 248748 393718
rect 248696 393654 248748 393660
rect 248708 16250 248736 393654
rect 248800 22982 248828 393858
rect 248788 22976 248840 22982
rect 248788 22918 248840 22924
rect 248892 22914 248920 393944
rect 249076 393802 249104 400044
rect 248984 393774 249104 393802
rect 248984 28286 249012 393774
rect 249168 393718 249196 400044
rect 249260 395690 249288 400044
rect 249248 395684 249300 395690
rect 249248 395626 249300 395632
rect 249248 395072 249300 395078
rect 249248 395014 249300 395020
rect 249156 393712 249208 393718
rect 249156 393654 249208 393660
rect 249260 391270 249288 395014
rect 249352 393786 249380 400044
rect 249340 393780 249392 393786
rect 249340 393722 249392 393728
rect 249248 391264 249300 391270
rect 249248 391206 249300 391212
rect 249444 389174 249472 400044
rect 249536 397633 249564 400044
rect 249522 397624 249578 397633
rect 249522 397559 249578 397568
rect 249628 397497 249656 400044
rect 249720 397769 249748 400044
rect 249706 397760 249762 397769
rect 249706 397695 249762 397704
rect 249614 397488 249670 397497
rect 249614 397423 249670 397432
rect 249812 393922 249840 400044
rect 249904 398041 249932 400044
rect 249890 398032 249946 398041
rect 249890 397967 249946 397976
rect 249892 394596 249944 394602
rect 249892 394538 249944 394544
rect 249800 393916 249852 393922
rect 249800 393858 249852 393864
rect 249904 393802 249932 394538
rect 249076 389146 249472 389174
rect 249812 393774 249932 393802
rect 249076 89010 249104 389146
rect 249064 89004 249116 89010
rect 249064 88946 249116 88952
rect 248972 28280 249024 28286
rect 248972 28222 249024 28228
rect 248880 22908 248932 22914
rect 248880 22850 248932 22856
rect 248696 16244 248748 16250
rect 248696 16186 248748 16192
rect 249812 16114 249840 393774
rect 249996 392442 250024 400044
rect 249904 392414 250024 392442
rect 249904 16182 249932 392414
rect 249984 392352 250036 392358
rect 249984 392294 250036 392300
rect 249892 16176 249944 16182
rect 249892 16118 249944 16124
rect 249800 16108 249852 16114
rect 249800 16050 249852 16056
rect 249996 16046 250024 392294
rect 250088 22778 250116 400044
rect 250180 394534 250208 400044
rect 250272 394602 250300 400044
rect 250364 395622 250392 400044
rect 250352 395616 250404 395622
rect 250352 395558 250404 395564
rect 250260 394596 250312 394602
rect 250260 394538 250312 394544
rect 250168 394528 250220 394534
rect 250168 394470 250220 394476
rect 250456 394210 250484 400044
rect 250364 394182 250484 394210
rect 250168 393916 250220 393922
rect 250168 393858 250220 393864
rect 250260 393916 250312 393922
rect 250260 393858 250312 393864
rect 250180 22846 250208 393858
rect 250272 24410 250300 393858
rect 250364 86290 250392 394182
rect 250548 392358 250576 400044
rect 250640 393922 250668 400044
rect 250628 393916 250680 393922
rect 250628 393858 250680 393864
rect 250536 392352 250588 392358
rect 250536 392294 250588 392300
rect 250732 392170 250760 400044
rect 250824 397497 250852 400044
rect 250916 397905 250944 400044
rect 250902 397896 250958 397905
rect 250902 397831 250958 397840
rect 251008 397769 251036 400044
rect 250994 397760 251050 397769
rect 250994 397695 251050 397704
rect 251100 397633 251128 400044
rect 251086 397624 251142 397633
rect 251086 397559 251142 397568
rect 250810 397488 250866 397497
rect 250810 397423 250866 397432
rect 250812 394528 250864 394534
rect 250812 394470 250864 394476
rect 250456 392142 250760 392170
rect 250456 177410 250484 392142
rect 250824 389174 250852 394470
rect 251192 392358 251220 400044
rect 251284 398313 251312 400044
rect 251270 398304 251326 398313
rect 251270 398239 251326 398248
rect 251272 398200 251324 398206
rect 251272 398142 251324 398148
rect 251284 397798 251312 398142
rect 251272 397792 251324 397798
rect 251272 397734 251324 397740
rect 251376 393972 251404 400044
rect 251468 395554 251496 400044
rect 251456 395548 251508 395554
rect 251456 395490 251508 395496
rect 251560 394670 251588 400044
rect 251548 394664 251600 394670
rect 251548 394606 251600 394612
rect 251548 394528 251600 394534
rect 251548 394470 251600 394476
rect 251376 393944 251496 393972
rect 251364 393848 251416 393854
rect 251364 393790 251416 393796
rect 251272 393780 251324 393786
rect 251272 393722 251324 393728
rect 251180 392352 251232 392358
rect 251180 392294 251232 392300
rect 250548 389146 250852 389174
rect 250548 352646 250576 389146
rect 250536 352640 250588 352646
rect 250536 352582 250588 352588
rect 250444 177404 250496 177410
rect 250444 177346 250496 177352
rect 250352 86284 250404 86290
rect 250352 86226 250404 86232
rect 250260 24404 250312 24410
rect 250260 24346 250312 24352
rect 250168 22840 250220 22846
rect 250168 22782 250220 22788
rect 250076 22772 250128 22778
rect 250076 22714 250128 22720
rect 249984 16040 250036 16046
rect 249984 15982 250036 15988
rect 248604 14544 248656 14550
rect 248604 14486 248656 14492
rect 248420 5092 248472 5098
rect 248420 5034 248472 5040
rect 251284 5030 251312 393722
rect 251376 15910 251404 393790
rect 251468 15978 251496 393944
rect 251560 17542 251588 394470
rect 251652 393854 251680 400044
rect 251744 393922 251772 400044
rect 251732 393916 251784 393922
rect 251732 393858 251784 393864
rect 251640 393848 251692 393854
rect 251640 393790 251692 393796
rect 251836 392442 251864 400044
rect 251928 394534 251956 400044
rect 252020 395486 252048 400044
rect 252008 395480 252060 395486
rect 252008 395422 252060 395428
rect 251916 394528 251968 394534
rect 251916 394470 251968 394476
rect 251916 393916 251968 393922
rect 251916 393858 251968 393864
rect 251744 392414 251864 392442
rect 251640 354000 251692 354006
rect 251640 353942 251692 353948
rect 251548 17536 251600 17542
rect 251548 17478 251600 17484
rect 251652 16574 251680 353942
rect 251744 177342 251772 392414
rect 251824 392352 251876 392358
rect 251824 392294 251876 392300
rect 251836 352578 251864 392294
rect 251928 354074 251956 393858
rect 252112 393786 252140 400044
rect 252204 397769 252232 400044
rect 252190 397760 252246 397769
rect 252190 397695 252246 397704
rect 252296 397633 252324 400044
rect 252282 397624 252338 397633
rect 252282 397559 252338 397568
rect 252388 397497 252416 400044
rect 252480 397905 252508 400044
rect 252466 397896 252522 397905
rect 252466 397831 252522 397840
rect 252374 397488 252430 397497
rect 252374 397423 252430 397432
rect 252192 394664 252244 394670
rect 252192 394606 252244 394612
rect 252100 393780 252152 393786
rect 252100 393722 252152 393728
rect 251916 354068 251968 354074
rect 251916 354010 251968 354016
rect 251824 352572 251876 352578
rect 251824 352514 251876 352520
rect 251732 177336 251784 177342
rect 251732 177278 251784 177284
rect 252204 16574 252232 394606
rect 252572 394074 252600 400044
rect 252664 399566 252692 400044
rect 252652 399560 252704 399566
rect 252652 399502 252704 399508
rect 252652 399424 252704 399430
rect 252652 399366 252704 399372
rect 252480 394046 252600 394074
rect 252480 393718 252508 394046
rect 252664 393972 252692 399366
rect 252572 393944 252692 393972
rect 252468 393712 252520 393718
rect 252468 393654 252520 393660
rect 251652 16546 252140 16574
rect 252204 16546 252508 16574
rect 251456 15972 251508 15978
rect 251456 15914 251508 15920
rect 251364 15904 251416 15910
rect 251364 15846 251416 15852
rect 251272 5024 251324 5030
rect 251272 4966 251324 4972
rect 248788 4888 248840 4894
rect 248788 4830 248840 4836
rect 248052 3528 248104 3534
rect 248052 3470 248104 3476
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247592 3392 247644 3398
rect 247592 3334 247644 3340
rect 247604 480 247632 3334
rect 248800 480 248828 4830
rect 251180 4820 251232 4826
rect 251180 4762 251232 4768
rect 249984 3052 250036 3058
rect 249984 2994 250036 3000
rect 249996 480 250024 2994
rect 251192 480 251220 4762
rect 252112 3482 252140 16546
rect 252112 3454 252416 3482
rect 252480 3466 252508 16546
rect 252572 4894 252600 393944
rect 252652 393848 252704 393854
rect 252652 393790 252704 393796
rect 252664 4962 252692 393790
rect 252756 17474 252784 400044
rect 252848 394534 252876 400044
rect 252836 394528 252888 394534
rect 252836 394470 252888 394476
rect 252940 394074 252968 400044
rect 252848 394046 252968 394074
rect 252848 393854 252876 394046
rect 253032 393972 253060 400044
rect 253124 399401 253152 400044
rect 253216 399430 253244 400044
rect 253204 399424 253256 399430
rect 253110 399392 253166 399401
rect 253204 399366 253256 399372
rect 253110 399327 253166 399336
rect 253112 399220 253164 399226
rect 253112 399162 253164 399168
rect 253204 399220 253256 399226
rect 253204 399162 253256 399168
rect 253124 398546 253152 399162
rect 253216 398818 253244 399162
rect 253204 398812 253256 398818
rect 253204 398754 253256 398760
rect 253202 398712 253258 398721
rect 253202 398647 253258 398656
rect 253112 398540 253164 398546
rect 253112 398482 253164 398488
rect 253110 398304 253166 398313
rect 253110 398239 253166 398248
rect 253124 397866 253152 398239
rect 253112 397860 253164 397866
rect 253112 397802 253164 397808
rect 253216 395418 253244 398647
rect 253204 395412 253256 395418
rect 253204 395354 253256 395360
rect 253204 394528 253256 394534
rect 253204 394470 253256 394476
rect 252940 393944 253060 393972
rect 252836 393848 252888 393854
rect 252836 393790 252888 393796
rect 252836 391060 252888 391066
rect 252836 391002 252888 391008
rect 252744 17468 252796 17474
rect 252744 17410 252796 17416
rect 252848 17338 252876 391002
rect 252940 17406 252968 393944
rect 253020 393848 253072 393854
rect 253020 393790 253072 393796
rect 253032 24206 253060 393790
rect 253112 393712 253164 393718
rect 253112 393654 253164 393660
rect 253124 24342 253152 393654
rect 253112 24336 253164 24342
rect 253112 24278 253164 24284
rect 253216 24274 253244 394470
rect 253308 391066 253336 400044
rect 253400 393854 253428 400044
rect 253388 393848 253440 393854
rect 253388 393790 253440 393796
rect 253296 391060 253348 391066
rect 253296 391002 253348 391008
rect 253492 389174 253520 400044
rect 253584 397497 253612 400044
rect 253676 399537 253704 400044
rect 253662 399528 253718 399537
rect 253662 399463 253718 399472
rect 253664 399356 253716 399362
rect 253664 399298 253716 399304
rect 253676 398682 253704 399298
rect 253664 398676 253716 398682
rect 253664 398618 253716 398624
rect 253662 398440 253718 398449
rect 253662 398375 253718 398384
rect 253676 397905 253704 398375
rect 253662 397896 253718 397905
rect 253662 397831 253718 397840
rect 253768 397769 253796 400044
rect 253754 397760 253810 397769
rect 253754 397695 253810 397704
rect 253860 397633 253888 400044
rect 253846 397624 253902 397633
rect 253846 397559 253902 397568
rect 253570 397488 253626 397497
rect 253570 397423 253626 397432
rect 253952 394806 253980 400044
rect 254044 398138 254072 400044
rect 254032 398132 254084 398138
rect 254032 398074 254084 398080
rect 254032 397928 254084 397934
rect 254032 397870 254084 397876
rect 254044 397730 254072 397870
rect 254032 397724 254084 397730
rect 254032 397666 254084 397672
rect 253940 394800 253992 394806
rect 253940 394742 253992 394748
rect 253940 394664 253992 394670
rect 254136 394618 254164 400044
rect 253940 394606 253992 394612
rect 253308 389146 253520 389174
rect 253308 351218 253336 389146
rect 253296 351212 253348 351218
rect 253296 351154 253348 351160
rect 253204 24268 253256 24274
rect 253204 24210 253256 24216
rect 253020 24200 253072 24206
rect 253020 24142 253072 24148
rect 252928 17400 252980 17406
rect 252928 17342 252980 17348
rect 252836 17332 252888 17338
rect 252836 17274 252888 17280
rect 253952 6254 253980 394606
rect 254044 394590 254164 394618
rect 254044 393718 254072 394590
rect 254124 394528 254176 394534
rect 254124 394470 254176 394476
rect 254032 393712 254084 393718
rect 254032 393654 254084 393660
rect 254032 393576 254084 393582
rect 254032 393518 254084 393524
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254044 6186 254072 393518
rect 254136 8974 254164 394470
rect 254228 393938 254256 400044
rect 254320 397594 254348 400044
rect 254308 397588 254360 397594
rect 254308 397530 254360 397536
rect 254412 394534 254440 400044
rect 254400 394528 254452 394534
rect 254400 394470 254452 394476
rect 254228 393910 254440 393938
rect 254308 393848 254360 393854
rect 254308 393790 254360 393796
rect 254216 393780 254268 393786
rect 254216 393722 254268 393728
rect 254228 14482 254256 393722
rect 254320 17270 254348 393790
rect 254412 24138 254440 393910
rect 254504 393854 254532 400044
rect 254596 394670 254624 400044
rect 254584 394664 254636 394670
rect 254584 394606 254636 394612
rect 254584 393916 254636 393922
rect 254584 393858 254636 393864
rect 254492 393848 254544 393854
rect 254492 393790 254544 393796
rect 254492 393712 254544 393718
rect 254492 393654 254544 393660
rect 254504 84862 254532 393654
rect 254596 347070 254624 393858
rect 254688 393786 254716 400044
rect 254780 399702 254808 400044
rect 254768 399696 254820 399702
rect 254768 399638 254820 399644
rect 254768 399560 254820 399566
rect 254768 399502 254820 399508
rect 254780 398206 254808 399502
rect 254768 398200 254820 398206
rect 254768 398142 254820 398148
rect 254768 394800 254820 394806
rect 254768 394742 254820 394748
rect 254676 393780 254728 393786
rect 254676 393722 254728 393728
rect 254780 389174 254808 394742
rect 254872 393582 254900 400044
rect 254964 393922 254992 400044
rect 255056 397497 255084 400044
rect 255148 397633 255176 400044
rect 255240 399265 255268 400044
rect 255226 399256 255282 399265
rect 255226 399191 255282 399200
rect 255228 398812 255280 398818
rect 255228 398754 255280 398760
rect 255134 397624 255190 397633
rect 255134 397559 255190 397568
rect 255042 397488 255098 397497
rect 255042 397423 255098 397432
rect 255240 395350 255268 398754
rect 255228 395344 255280 395350
rect 255228 395286 255280 395292
rect 255332 393938 255360 400044
rect 255424 398410 255452 400044
rect 255412 398404 255464 398410
rect 255412 398346 255464 398352
rect 254952 393916 255004 393922
rect 255332 393910 255452 393938
rect 254952 393858 255004 393864
rect 255320 393848 255372 393854
rect 255320 393790 255372 393796
rect 254860 393576 254912 393582
rect 254860 393518 254912 393524
rect 254688 389146 254808 389174
rect 254688 354006 254716 389146
rect 254676 354000 254728 354006
rect 254676 353942 254728 353948
rect 254584 347064 254636 347070
rect 254584 347006 254636 347012
rect 254492 84856 254544 84862
rect 254492 84798 254544 84804
rect 254400 24132 254452 24138
rect 254400 24074 254452 24080
rect 254308 17264 254360 17270
rect 254308 17206 254360 17212
rect 254216 14476 254268 14482
rect 254216 14418 254268 14424
rect 254124 8968 254176 8974
rect 254124 8910 254176 8916
rect 254032 6180 254084 6186
rect 254032 6122 254084 6128
rect 254674 5400 254730 5409
rect 254674 5335 254730 5344
rect 252652 4956 252704 4962
rect 252652 4898 252704 4904
rect 252560 4888 252612 4894
rect 252560 4830 252612 4836
rect 253480 3596 253532 3602
rect 253480 3538 253532 3544
rect 252388 480 252416 3454
rect 252468 3460 252520 3466
rect 252468 3402 252520 3408
rect 253492 480 253520 3538
rect 254688 480 254716 5335
rect 255332 3482 255360 393790
rect 255424 4826 255452 393910
rect 255516 10334 255544 400044
rect 255608 398313 255636 400044
rect 255688 399696 255740 399702
rect 255688 399638 255740 399644
rect 255700 398818 255728 399638
rect 257250 399120 257306 399129
rect 257250 399055 257306 399064
rect 255688 398812 255740 398818
rect 255688 398754 255740 398760
rect 257264 398721 257292 399055
rect 257712 398744 257764 398750
rect 257250 398712 257306 398721
rect 256056 398676 256108 398682
rect 257712 398686 257764 398692
rect 257250 398647 257306 398656
rect 256056 398618 256108 398624
rect 255594 398304 255650 398313
rect 255594 398239 255650 398248
rect 255594 395720 255650 395729
rect 255594 395655 255650 395664
rect 255608 393854 255636 395655
rect 255964 394596 256016 394602
rect 255964 394538 256016 394544
rect 255596 393848 255648 393854
rect 255596 393790 255648 393796
rect 255504 10328 255556 10334
rect 255504 10270 255556 10276
rect 255412 4820 255464 4826
rect 255412 4762 255464 4768
rect 255976 3602 256004 394538
rect 256068 26926 256096 398618
rect 256238 398576 256294 398585
rect 256238 398511 256294 398520
rect 256148 398064 256200 398070
rect 256148 398006 256200 398012
rect 256160 26994 256188 398006
rect 256252 28354 256280 398511
rect 256700 398336 256752 398342
rect 256700 398278 256752 398284
rect 256790 398304 256846 398313
rect 256240 28348 256292 28354
rect 256240 28290 256292 28296
rect 256148 26988 256200 26994
rect 256148 26930 256200 26936
rect 256056 26920 256108 26926
rect 256056 26862 256108 26868
rect 255964 3596 256016 3602
rect 255964 3538 256016 3544
rect 255332 3454 255912 3482
rect 255884 480 255912 3454
rect 256712 3058 256740 398278
rect 256790 398239 256846 398248
rect 257528 398268 257580 398274
rect 256804 397526 256832 398239
rect 257528 398210 257580 398216
rect 257436 397656 257488 397662
rect 257436 397598 257488 397604
rect 256792 397520 256844 397526
rect 256792 397462 256844 397468
rect 257344 397316 257396 397322
rect 257344 397258 257396 397264
rect 257356 3670 257384 397258
rect 257448 7682 257476 397598
rect 257436 7676 257488 7682
rect 257436 7618 257488 7624
rect 257540 7614 257568 398210
rect 257620 392896 257672 392902
rect 257620 392838 257672 392844
rect 257528 7608 257580 7614
rect 257528 7550 257580 7556
rect 257632 3874 257660 392838
rect 257724 352714 257752 398686
rect 258814 398576 258870 398585
rect 258814 398511 258870 398520
rect 258724 397724 258776 397730
rect 258724 397666 258776 397672
rect 257712 352708 257764 352714
rect 257712 352650 257764 352656
rect 258736 35222 258764 397666
rect 258828 302938 258856 398511
rect 260024 398342 260052 400143
rect 263506 398712 263562 398721
rect 263506 398647 263562 398656
rect 262864 398472 262916 398478
rect 262864 398414 262916 398420
rect 263414 398440 263470 398449
rect 260012 398336 260064 398342
rect 260012 398278 260064 398284
rect 260196 397996 260248 398002
rect 260196 397938 260248 397944
rect 260104 397928 260156 397934
rect 260104 397870 260156 397876
rect 259460 397792 259512 397798
rect 259460 397734 259512 397740
rect 258816 302932 258868 302938
rect 258816 302874 258868 302880
rect 258724 35216 258776 35222
rect 258724 35158 258776 35164
rect 259472 11694 259500 397734
rect 259552 352844 259604 352850
rect 259552 352786 259604 352792
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 352786
rect 260116 49026 260144 397870
rect 260208 336054 260236 397938
rect 261482 397760 261538 397769
rect 261482 397695 261538 397704
rect 260196 336048 260248 336054
rect 260196 335990 260248 335996
rect 260104 49020 260156 49026
rect 260104 48962 260156 48968
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 258262 5264 258318 5273
rect 258262 5199 258318 5208
rect 257620 3868 257672 3874
rect 257620 3810 257672 3816
rect 257068 3664 257120 3670
rect 257068 3606 257120 3612
rect 257344 3664 257396 3670
rect 257344 3606 257396 3612
rect 256700 3052 256752 3058
rect 256700 2994 256752 3000
rect 257080 480 257108 3606
rect 258276 480 258304 5199
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261496 9042 261524 397695
rect 262876 182850 262904 398414
rect 263520 398426 263548 398647
rect 263470 398398 263548 398426
rect 263414 398375 263470 398384
rect 262864 182844 262916 182850
rect 262864 182786 262916 182792
rect 264256 86970 264284 444751
rect 264336 443216 264388 443222
rect 264336 443158 264388 443164
rect 264348 206990 264376 443158
rect 264440 399090 264468 446247
rect 264532 399158 264560 446694
rect 264612 443488 264664 443494
rect 264612 443430 264664 443436
rect 264624 401266 264652 443430
rect 264612 401260 264664 401266
rect 264612 401202 264664 401208
rect 264716 400994 264744 446762
rect 265806 445904 265862 445913
rect 265806 445839 265862 445848
rect 265714 444680 265770 444689
rect 265714 444615 265770 444624
rect 265256 443624 265308 443630
rect 265256 443566 265308 443572
rect 265622 443592 265678 443601
rect 265268 436082 265296 443566
rect 265622 443527 265678 443536
rect 265256 436076 265308 436082
rect 265256 436018 265308 436024
rect 264704 400988 264756 400994
rect 264704 400930 264756 400936
rect 264520 399152 264572 399158
rect 264520 399094 264572 399100
rect 264428 399084 264480 399090
rect 264428 399026 264480 399032
rect 264336 206984 264388 206990
rect 264336 206926 264388 206932
rect 264244 86964 264296 86970
rect 264244 86906 264296 86912
rect 262220 82204 262272 82210
rect 262220 82146 262272 82152
rect 262232 16574 262260 82146
rect 265636 73166 265664 443527
rect 265728 113150 265756 444615
rect 265820 233238 265848 445839
rect 265912 400926 265940 446830
rect 267002 444544 267058 444553
rect 267002 444479 267058 444488
rect 265992 444440 266044 444446
rect 265992 444382 266044 444388
rect 266004 431934 266032 444382
rect 265992 431928 266044 431934
rect 265992 431870 266044 431876
rect 265900 400920 265952 400926
rect 265900 400862 265952 400868
rect 266360 352776 266412 352782
rect 266360 352718 266412 352724
rect 265808 233232 265860 233238
rect 265808 233174 265860 233180
rect 265716 113144 265768 113150
rect 265716 113086 265768 113092
rect 265624 73160 265676 73166
rect 265624 73102 265676 73108
rect 266372 16574 266400 352718
rect 267016 126954 267044 444479
rect 267108 398750 267136 448462
rect 281644 446554 281672 591194
rect 281736 446622 281764 596838
rect 281814 596799 281870 596808
rect 281828 449342 281856 596799
rect 281816 449336 281868 449342
rect 281816 449278 281868 449284
rect 281920 449002 281948 596974
rect 282000 596964 282052 596970
rect 282000 596906 282052 596912
rect 282012 596358 282040 596906
rect 282104 596358 282132 597110
rect 282196 596834 282224 597178
rect 282276 596896 282328 596902
rect 282276 596838 282328 596844
rect 282184 596828 282236 596834
rect 282184 596770 282236 596776
rect 282000 596352 282052 596358
rect 282000 596294 282052 596300
rect 282092 596352 282144 596358
rect 282092 596294 282144 596300
rect 282000 591388 282052 591394
rect 282000 591330 282052 591336
rect 282012 449818 282040 591330
rect 282000 449812 282052 449818
rect 282000 449754 282052 449760
rect 282104 449070 282132 596294
rect 282196 449682 282224 596770
rect 282288 596426 282316 596838
rect 282276 596420 282328 596426
rect 282276 596362 282328 596368
rect 282184 449676 282236 449682
rect 282184 449618 282236 449624
rect 282288 449546 282316 596362
rect 282380 591258 282408 597518
rect 284666 597272 284722 597281
rect 284666 597207 284722 597216
rect 284300 597100 284352 597106
rect 284300 597042 284352 597048
rect 284312 596562 284340 597042
rect 284390 597000 284446 597009
rect 284680 596970 284708 597207
rect 284758 597136 284814 597145
rect 284758 597071 284814 597080
rect 284390 596935 284446 596944
rect 284668 596964 284720 596970
rect 284300 596556 284352 596562
rect 284300 596498 284352 596504
rect 282368 591252 282420 591258
rect 282368 591194 282420 591200
rect 283564 590708 283616 590714
rect 283564 590650 283616 590656
rect 282828 518220 282880 518226
rect 282828 518162 282880 518168
rect 282840 489914 282868 518162
rect 282380 489886 282868 489914
rect 282380 488073 282408 489886
rect 282366 488064 282422 488073
rect 282366 487999 282422 488008
rect 282380 478242 282408 487999
rect 282368 478236 282420 478242
rect 282368 478178 282420 478184
rect 283576 453558 283604 590650
rect 284208 523728 284260 523734
rect 284208 523670 284260 523676
rect 284116 521008 284168 521014
rect 284116 520950 284168 520956
rect 284024 520940 284076 520946
rect 284024 520882 284076 520888
rect 284036 489802 284064 520882
rect 284024 489796 284076 489802
rect 284024 489738 284076 489744
rect 283656 488708 283708 488714
rect 283656 488650 283708 488656
rect 283564 453552 283616 453558
rect 283564 453494 283616 453500
rect 283668 451246 283696 488650
rect 284036 479602 284064 489738
rect 284128 489734 284156 520950
rect 284220 489802 284248 523670
rect 284208 489796 284260 489802
rect 284208 489738 284260 489744
rect 284116 489728 284168 489734
rect 284116 489670 284168 489676
rect 284128 481030 284156 489670
rect 284220 488714 284248 489738
rect 284208 488708 284260 488714
rect 284208 488650 284260 488656
rect 284116 481024 284168 481030
rect 284116 480966 284168 480972
rect 284024 479596 284076 479602
rect 284024 479538 284076 479544
rect 283656 451240 283708 451246
rect 283656 451182 283708 451188
rect 284312 449750 284340 596498
rect 284404 596494 284432 596935
rect 284668 596906 284720 596912
rect 284576 596692 284628 596698
rect 284576 596634 284628 596640
rect 284484 596624 284536 596630
rect 284484 596566 284536 596572
rect 284392 596488 284444 596494
rect 284392 596430 284444 596436
rect 284300 449744 284352 449750
rect 284300 449686 284352 449692
rect 282276 449540 282328 449546
rect 282276 449482 282328 449488
rect 284404 449410 284432 596430
rect 284496 449886 284524 596566
rect 284588 596562 284616 596634
rect 284576 596556 284628 596562
rect 284576 596498 284628 596504
rect 284484 449880 284536 449886
rect 284484 449822 284536 449828
rect 284392 449404 284444 449410
rect 284392 449346 284444 449352
rect 284588 449138 284616 596498
rect 284680 449313 284708 596906
rect 284772 596290 284800 597071
rect 284944 596828 284996 596834
rect 284944 596770 284996 596776
rect 284760 596284 284812 596290
rect 284760 596226 284812 596232
rect 284666 449304 284722 449313
rect 284666 449239 284722 449248
rect 284772 449177 284800 596226
rect 284956 596222 284984 596770
rect 284944 596216 284996 596222
rect 284944 596158 284996 596164
rect 284956 586514 284984 596158
rect 284864 586486 284984 586514
rect 284864 449614 284892 586486
rect 284944 526448 284996 526454
rect 284944 526390 284996 526396
rect 284956 484362 284984 526390
rect 285588 523796 285640 523802
rect 285588 523738 285640 523744
rect 285600 489841 285628 523738
rect 285586 489832 285642 489841
rect 285586 489767 285642 489776
rect 285600 488617 285628 489767
rect 285034 488608 285090 488617
rect 285034 488543 285090 488552
rect 285586 488608 285642 488617
rect 285586 488543 285642 488552
rect 284944 484356 284996 484362
rect 284944 484298 284996 484304
rect 285048 452606 285076 488543
rect 290476 454850 290504 696934
rect 290568 472666 290596 700334
rect 294604 700324 294656 700330
rect 294604 700266 294656 700272
rect 290556 472660 290608 472666
rect 290556 472602 290608 472608
rect 290464 454844 290516 454850
rect 290464 454786 290516 454792
rect 285036 452600 285088 452606
rect 285036 452542 285088 452548
rect 294616 450702 294644 700266
rect 298744 699712 298796 699718
rect 298744 699654 298796 699660
rect 298006 636984 298062 636993
rect 298006 636919 298062 636928
rect 297914 635896 297970 635905
rect 297914 635831 297970 635840
rect 297822 634264 297878 634273
rect 297822 634199 297878 634208
rect 297638 633176 297694 633185
rect 297638 633111 297694 633120
rect 297454 631544 297510 631553
rect 297454 631479 297510 631488
rect 296994 610192 297050 610201
rect 296994 610127 297050 610136
rect 296902 608288 296958 608297
rect 296902 608223 296958 608232
rect 294696 525972 294748 525978
rect 294696 525914 294748 525920
rect 294708 482390 294736 525914
rect 296916 498273 296944 608223
rect 297008 500857 297036 610127
rect 297086 608696 297142 608705
rect 297086 608631 297142 608640
rect 296994 500848 297050 500857
rect 296994 500783 297050 500792
rect 297100 499574 297128 608631
rect 297364 599820 297416 599826
rect 297364 599762 297416 599768
rect 297272 599412 297324 599418
rect 297272 599354 297324 599360
rect 297180 598324 297232 598330
rect 297180 598266 297232 598272
rect 297192 526454 297220 598266
rect 297180 526448 297232 526454
rect 297180 526390 297232 526396
rect 297284 525978 297312 599354
rect 297272 525972 297324 525978
rect 297272 525914 297324 525920
rect 297376 523802 297404 599762
rect 297468 598942 297496 631479
rect 297546 628552 297602 628561
rect 297546 628487 297602 628496
rect 297456 598936 297508 598942
rect 297456 598878 297508 598884
rect 297364 523796 297416 523802
rect 297364 523738 297416 523744
rect 297468 521665 297496 598878
rect 297560 598874 297588 628487
rect 297548 598868 297600 598874
rect 297548 598810 297600 598816
rect 297454 521656 297510 521665
rect 297454 521591 297510 521600
rect 297468 521014 297496 521591
rect 297456 521008 297508 521014
rect 297456 520950 297508 520956
rect 297560 518673 297588 598810
rect 297652 523734 297680 633111
rect 297730 630184 297786 630193
rect 297730 630119 297786 630128
rect 297744 538214 297772 630119
rect 297836 600030 297864 634199
rect 297824 600024 297876 600030
rect 297824 599966 297876 599972
rect 297836 599826 297864 599966
rect 297824 599820 297876 599826
rect 297824 599762 297876 599768
rect 297928 599622 297956 635831
rect 297916 599616 297968 599622
rect 297916 599558 297968 599564
rect 297928 599418 297956 599558
rect 297916 599412 297968 599418
rect 297916 599354 297968 599360
rect 298020 598330 298048 636919
rect 298008 598324 298060 598330
rect 298008 598266 298060 598272
rect 297744 538186 297864 538214
rect 297730 527096 297786 527105
rect 297730 527031 297786 527040
rect 297744 526454 297772 527031
rect 297732 526448 297784 526454
rect 297732 526390 297784 526396
rect 297640 523728 297692 523734
rect 297640 523670 297692 523676
rect 297836 520946 297864 538186
rect 298006 526008 298062 526017
rect 298006 525943 298008 525952
rect 298060 525943 298062 525952
rect 298008 525914 298060 525920
rect 298006 524376 298062 524385
rect 298006 524311 298062 524320
rect 298020 523802 298048 524311
rect 298008 523796 298060 523802
rect 298008 523738 298060 523744
rect 297916 523728 297968 523734
rect 297916 523670 297968 523676
rect 297928 523297 297956 523670
rect 297914 523288 297970 523297
rect 297914 523223 297970 523232
rect 297824 520940 297876 520946
rect 297824 520882 297876 520888
rect 297836 520305 297864 520882
rect 297822 520296 297878 520305
rect 297822 520231 297878 520240
rect 297546 518664 297602 518673
rect 297546 518599 297602 518608
rect 297560 518226 297588 518599
rect 297548 518220 297600 518226
rect 297548 518162 297600 518168
rect 297914 500848 297970 500857
rect 297914 500783 297970 500792
rect 297928 500313 297956 500783
rect 297914 500304 297970 500313
rect 297914 500239 297970 500248
rect 297100 499546 297496 499574
rect 297468 498681 297496 499546
rect 297454 498672 297510 498681
rect 297454 498607 297510 498616
rect 296902 498264 296958 498273
rect 296902 498199 296958 498208
rect 297364 488708 297416 488714
rect 297364 488650 297416 488656
rect 294696 482384 294748 482390
rect 294696 482326 294748 482332
rect 295984 458720 296036 458726
rect 295984 458662 296036 458668
rect 294604 450696 294656 450702
rect 294604 450638 294656 450644
rect 284852 449608 284904 449614
rect 284852 449550 284904 449556
rect 284758 449168 284814 449177
rect 284576 449132 284628 449138
rect 284758 449103 284814 449112
rect 284576 449074 284628 449080
rect 282092 449064 282144 449070
rect 282092 449006 282144 449012
rect 281908 448996 281960 449002
rect 281908 448938 281960 448944
rect 295996 447846 296024 458662
rect 297376 448526 297404 488650
rect 297468 480962 297496 498607
rect 297822 498264 297878 498273
rect 297822 498199 297878 498208
rect 297836 489598 297864 498199
rect 297928 489666 297956 500239
rect 297916 489660 297968 489666
rect 297916 489602 297968 489608
rect 297824 489592 297876 489598
rect 297824 489534 297876 489540
rect 297836 488714 297864 489534
rect 297824 488708 297876 488714
rect 297824 488650 297876 488656
rect 297928 485110 297956 489602
rect 297916 485104 297968 485110
rect 297916 485046 297968 485052
rect 297456 480956 297508 480962
rect 297456 480898 297508 480904
rect 298652 476060 298704 476066
rect 298652 476002 298704 476008
rect 298664 475454 298692 476002
rect 298652 475448 298704 475454
rect 298652 475390 298704 475396
rect 298652 471980 298704 471986
rect 298652 471922 298704 471928
rect 298664 471306 298692 471922
rect 298652 471300 298704 471306
rect 298652 471242 298704 471248
rect 297548 458448 297600 458454
rect 297548 458390 297600 458396
rect 297560 453354 297588 458390
rect 298756 453490 298784 699654
rect 298848 467294 298876 700402
rect 300136 699718 300164 703520
rect 332520 700466 332548 703520
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364996 700330 365024 703520
rect 392584 700392 392636 700398
rect 392584 700334 392636 700340
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 335360 597576 335412 597582
rect 319994 597544 320050 597553
rect 319994 597479 320050 597488
rect 322294 597544 322350 597553
rect 322294 597479 322350 597488
rect 323398 597544 323454 597553
rect 323398 597479 323454 597488
rect 324778 597544 324834 597553
rect 324778 597479 324834 597488
rect 326158 597544 326214 597553
rect 326158 597479 326160 597488
rect 314658 597408 314714 597417
rect 314658 597343 314714 597352
rect 314672 596970 314700 597343
rect 299388 596964 299440 596970
rect 299388 596906 299440 596912
rect 314660 596964 314712 596970
rect 314660 596906 314712 596912
rect 299296 596284 299348 596290
rect 299296 596226 299348 596232
rect 299204 596216 299256 596222
rect 299204 596158 299256 596164
rect 299112 476468 299164 476474
rect 299112 476410 299164 476416
rect 299124 471986 299152 476410
rect 299216 476066 299244 596158
rect 299308 476354 299336 596226
rect 299400 476474 299428 596906
rect 320008 596902 320036 597479
rect 319996 596896 320048 596902
rect 319996 596838 320048 596844
rect 322308 596834 322336 597479
rect 323412 597174 323440 597479
rect 323400 597168 323452 597174
rect 323400 597110 323452 597116
rect 324792 597106 324820 597479
rect 326212 597479 326214 597488
rect 330390 597544 330446 597553
rect 330390 597479 330446 597488
rect 335358 597544 335360 597553
rect 335412 597544 335414 597553
rect 335358 597479 335414 597488
rect 340510 597544 340566 597553
rect 340510 597479 340566 597488
rect 345662 597544 345718 597553
rect 345662 597479 345718 597488
rect 350446 597544 350502 597553
rect 350446 597479 350502 597488
rect 354678 597544 354734 597553
rect 354678 597479 354734 597488
rect 360566 597544 360622 597553
rect 360566 597479 360622 597488
rect 326160 597450 326212 597456
rect 324320 597100 324372 597106
rect 324320 597042 324372 597048
rect 324780 597100 324832 597106
rect 324780 597042 324832 597048
rect 322296 596828 322348 596834
rect 322296 596770 322348 596776
rect 324332 596630 324360 597042
rect 324320 596624 324372 596630
rect 324320 596566 324372 596572
rect 326172 596562 326200 597450
rect 330404 597378 330432 597479
rect 330392 597372 330444 597378
rect 330392 597314 330444 597320
rect 330404 596766 330432 597314
rect 340524 597242 340552 597479
rect 345676 597310 345704 597479
rect 350460 597446 350488 597479
rect 350448 597440 350500 597446
rect 350448 597382 350500 597388
rect 345664 597304 345716 597310
rect 345664 597246 345716 597252
rect 340512 597236 340564 597242
rect 340512 597178 340564 597184
rect 354692 596766 354720 597479
rect 360580 597038 360608 597479
rect 360568 597032 360620 597038
rect 360568 596974 360620 596980
rect 330392 596760 330444 596766
rect 330392 596702 330444 596708
rect 354680 596760 354732 596766
rect 354680 596702 354732 596708
rect 326160 596556 326212 596562
rect 326160 596498 326212 596504
rect 311898 596320 311954 596329
rect 311898 596255 311900 596264
rect 311952 596255 311954 596264
rect 313278 596320 313334 596329
rect 313278 596255 313334 596264
rect 311900 596226 311952 596232
rect 313292 596222 313320 596255
rect 313280 596216 313332 596222
rect 313280 596158 313332 596164
rect 325330 489152 325386 489161
rect 325330 489087 325386 489096
rect 325344 488782 325372 489087
rect 325332 488776 325384 488782
rect 325332 488718 325384 488724
rect 336648 488776 336700 488782
rect 336648 488718 336700 488724
rect 336660 488646 336688 488718
rect 335452 488640 335504 488646
rect 335452 488582 335504 488588
rect 336648 488640 336700 488646
rect 336648 488582 336700 488588
rect 340604 488640 340656 488646
rect 340604 488582 340656 488588
rect 330484 488572 330536 488578
rect 330484 488514 330536 488520
rect 330496 488481 330524 488514
rect 335464 488481 335492 488582
rect 340616 488510 340644 488582
rect 340604 488504 340656 488510
rect 330482 488472 330538 488481
rect 330482 488407 330538 488416
rect 335450 488472 335506 488481
rect 335450 488407 335506 488416
rect 340602 488472 340604 488481
rect 340656 488472 340658 488481
rect 340602 488407 340658 488416
rect 345754 488472 345810 488481
rect 345754 488407 345810 488416
rect 350354 488472 350410 488481
rect 350354 488407 350410 488416
rect 355782 488472 355838 488481
rect 355782 488407 355838 488416
rect 360474 488472 360530 488481
rect 360474 488407 360530 488416
rect 313922 488336 313978 488345
rect 313922 488271 313978 488280
rect 312544 488232 312596 488238
rect 312544 488174 312596 488180
rect 312556 487257 312584 488174
rect 312542 487248 312598 487257
rect 312542 487183 312598 487192
rect 299388 476468 299440 476474
rect 299388 476410 299440 476416
rect 299308 476326 299428 476354
rect 299204 476060 299256 476066
rect 299204 476002 299256 476008
rect 299400 474638 299428 476326
rect 312556 474638 312584 487183
rect 313936 476066 313964 488271
rect 315302 488200 315358 488209
rect 315302 488135 315358 488144
rect 318892 488164 318944 488170
rect 313924 476060 313976 476066
rect 313924 476002 313976 476008
rect 299388 474632 299440 474638
rect 299388 474574 299440 474580
rect 312544 474632 312596 474638
rect 312544 474574 312596 474580
rect 299400 474026 299428 474574
rect 299388 474020 299440 474026
rect 299388 473962 299440 473968
rect 315316 471986 315344 488135
rect 318892 488106 318944 488112
rect 318904 487937 318932 488106
rect 326344 488096 326396 488102
rect 326344 488038 326396 488044
rect 318890 487928 318946 487937
rect 318890 487863 318946 487872
rect 318064 487756 318116 487762
rect 318064 487698 318116 487704
rect 318076 487257 318104 487698
rect 318062 487248 318118 487257
rect 318062 487183 318118 487192
rect 318076 473346 318104 487183
rect 318904 486470 318932 487863
rect 320824 487688 320876 487694
rect 320824 487630 320876 487636
rect 320088 487620 320140 487626
rect 320088 487562 320140 487568
rect 320100 487257 320128 487562
rect 320836 487257 320864 487630
rect 322204 487552 322256 487558
rect 322204 487494 322256 487500
rect 322216 487257 322244 487494
rect 323582 487384 323638 487393
rect 323582 487319 323638 487328
rect 323596 487286 323624 487319
rect 323584 487280 323636 487286
rect 319442 487248 319498 487257
rect 319442 487183 319498 487192
rect 320086 487248 320142 487257
rect 320086 487183 320142 487192
rect 320822 487248 320878 487257
rect 320822 487183 320878 487192
rect 322202 487248 322258 487257
rect 326356 487257 326384 488038
rect 345768 487966 345796 488407
rect 345756 487960 345808 487966
rect 345756 487902 345808 487908
rect 345768 487490 345796 487902
rect 350368 487830 350396 488407
rect 355796 487898 355824 488407
rect 360488 488034 360516 488407
rect 360476 488028 360528 488034
rect 360476 487970 360528 487976
rect 355784 487892 355836 487898
rect 355784 487834 355836 487840
rect 350356 487824 350408 487830
rect 350356 487766 350408 487772
rect 345756 487484 345808 487490
rect 345756 487426 345808 487432
rect 355796 487354 355824 487834
rect 360488 487422 360516 487970
rect 360476 487416 360528 487422
rect 360476 487358 360528 487364
rect 355784 487348 355836 487354
rect 355784 487290 355836 487296
rect 323584 487222 323636 487228
rect 324870 487248 324926 487257
rect 322202 487183 322258 487192
rect 318892 486464 318944 486470
rect 318892 486406 318944 486412
rect 319456 478854 319484 487183
rect 319444 478848 319496 478854
rect 319444 478790 319496 478796
rect 320836 474706 320864 487183
rect 322216 475386 322244 487183
rect 323596 476814 323624 487222
rect 324320 487212 324372 487218
rect 324870 487183 324872 487192
rect 324320 487154 324372 487160
rect 324924 487183 324926 487192
rect 326342 487248 326398 487257
rect 326342 487183 326398 487192
rect 324872 487154 324924 487160
rect 324332 482322 324360 487154
rect 324320 482316 324372 482322
rect 324320 482258 324372 482264
rect 326356 479534 326384 487183
rect 326344 479528 326396 479534
rect 326344 479470 326396 479476
rect 323584 476808 323636 476814
rect 323584 476750 323636 476756
rect 322204 475380 322256 475386
rect 322204 475322 322256 475328
rect 320824 474700 320876 474706
rect 320824 474642 320876 474648
rect 318064 473340 318116 473346
rect 318064 473282 318116 473288
rect 299112 471980 299164 471986
rect 299112 471922 299164 471928
rect 315304 471980 315356 471986
rect 315304 471922 315356 471928
rect 392596 469946 392624 700334
rect 393964 700324 394016 700330
rect 393964 700266 394016 700272
rect 392584 469940 392636 469946
rect 392584 469882 392636 469888
rect 298836 467288 298888 467294
rect 298836 467230 298888 467236
rect 393976 461854 394004 700266
rect 397472 465798 397500 703520
rect 402244 700528 402296 700534
rect 402244 700470 402296 700476
rect 397460 465792 397512 465798
rect 397460 465734 397512 465740
rect 402256 463078 402284 700470
rect 402336 700460 402388 700466
rect 402336 700402 402388 700408
rect 402348 469878 402376 700402
rect 413664 699718 413692 703520
rect 429856 700534 429884 703520
rect 429844 700528 429896 700534
rect 429844 700470 429896 700476
rect 462332 700466 462360 703520
rect 462320 700460 462372 700466
rect 462320 700402 462372 700408
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 505744 700324 505796 700330
rect 505744 700266 505796 700272
rect 409144 699712 409196 699718
rect 409144 699654 409196 699660
rect 413652 699712 413704 699718
rect 413652 699654 413704 699660
rect 407762 636440 407818 636449
rect 407762 636375 407818 636384
rect 407578 631000 407634 631009
rect 407578 630935 407634 630944
rect 407394 628008 407450 628017
rect 407394 627943 407450 627952
rect 407408 598874 407436 627943
rect 407592 598942 407620 630935
rect 407776 605834 407804 636375
rect 407946 635352 408002 635361
rect 407946 635287 408002 635296
rect 407854 607744 407910 607753
rect 407854 607679 407910 607688
rect 407684 605806 407804 605834
rect 407580 598936 407632 598942
rect 407580 598878 407632 598884
rect 407396 598868 407448 598874
rect 407396 598810 407448 598816
rect 407684 598754 407712 605806
rect 407764 600296 407816 600302
rect 407764 600238 407816 600244
rect 407776 599622 407804 600238
rect 407764 599616 407816 599622
rect 407764 599558 407816 599564
rect 407500 598726 407712 598754
rect 407500 598262 407528 598726
rect 407776 598618 407804 599558
rect 407684 598590 407804 598618
rect 407488 598256 407540 598262
rect 407488 598198 407540 598204
rect 407500 527105 407528 598198
rect 407486 527096 407542 527105
rect 407486 527031 407542 527040
rect 407684 526561 407712 598590
rect 407764 596216 407816 596222
rect 407764 596158 407816 596164
rect 407670 526552 407726 526561
rect 407670 526487 407726 526496
rect 407670 523288 407726 523297
rect 407670 523223 407726 523232
rect 407578 520976 407634 520985
rect 407578 520911 407634 520920
rect 407486 517984 407542 517993
rect 407486 517919 407542 517928
rect 407500 488073 407528 517919
rect 407592 489734 407620 520911
rect 407684 489802 407712 523223
rect 407672 489796 407724 489802
rect 407672 489738 407724 489744
rect 407580 489728 407632 489734
rect 407580 489670 407632 489676
rect 407776 488209 407804 596158
rect 407868 498409 407896 607679
rect 407960 600302 407988 635287
rect 408222 633720 408278 633729
rect 408222 633655 408278 633664
rect 408038 632632 408094 632641
rect 408038 632567 408094 632576
rect 407948 600296 408000 600302
rect 407948 600238 408000 600244
rect 407948 596284 408000 596290
rect 407948 596226 408000 596232
rect 407854 498400 407910 498409
rect 407854 498335 407910 498344
rect 407868 489598 407896 498335
rect 407856 489592 407908 489598
rect 407856 489534 407908 489540
rect 407960 488510 407988 596226
rect 408052 523297 408080 632567
rect 408130 629640 408186 629649
rect 408130 629575 408186 629584
rect 408038 523288 408094 523297
rect 408038 523223 408094 523232
rect 408144 520305 408172 629575
rect 408236 600030 408264 633655
rect 408406 610056 408462 610065
rect 408406 609991 408462 610000
rect 408314 608696 408370 608705
rect 408314 608631 408370 608640
rect 408224 600024 408276 600030
rect 408224 599966 408276 599972
rect 408224 596352 408276 596358
rect 408224 596294 408276 596300
rect 408130 520296 408186 520305
rect 408130 520231 408186 520240
rect 408038 498264 408094 498273
rect 408038 498199 408094 498208
rect 407948 488504 408000 488510
rect 407948 488446 408000 488452
rect 407960 488345 407988 488446
rect 407946 488336 408002 488345
rect 407946 488271 408002 488280
rect 407762 488200 407818 488209
rect 407762 488135 407818 488144
rect 407486 488064 407542 488073
rect 407486 487999 407542 488008
rect 402336 469872 402388 469878
rect 402336 469814 402388 469820
rect 408052 463146 408080 498199
rect 408144 489870 408172 520231
rect 408132 489864 408184 489870
rect 408132 489806 408184 489812
rect 408236 488442 408264 596294
rect 408328 498681 408356 608631
rect 408420 500313 408448 609991
rect 408406 500304 408462 500313
rect 408406 500239 408462 500248
rect 408314 498672 408370 498681
rect 408314 498607 408370 498616
rect 408328 498273 408356 498607
rect 408314 498264 408370 498273
rect 408314 498199 408370 498208
rect 408420 489666 408448 500239
rect 408408 489660 408460 489666
rect 408408 489602 408460 489608
rect 408224 488436 408276 488442
rect 408224 488378 408276 488384
rect 408236 488238 408264 488378
rect 408224 488232 408276 488238
rect 408224 488174 408276 488180
rect 409156 464506 409184 699654
rect 502984 670744 503036 670750
rect 502984 670686 503036 670692
rect 444380 597576 444432 597582
rect 429198 597544 429254 597553
rect 429198 597479 429254 597488
rect 434718 597544 434774 597553
rect 434718 597479 434720 597488
rect 429212 596902 429240 597479
rect 434772 597479 434774 597488
rect 444378 597544 444380 597553
rect 444432 597544 444434 597553
rect 444378 597479 444434 597488
rect 459558 597544 459614 597553
rect 459558 597479 459614 597488
rect 434720 597450 434772 597456
rect 459572 597446 459600 597479
rect 459560 597440 459612 597446
rect 440238 597408 440294 597417
rect 440238 597343 440240 597352
rect 440292 597343 440294 597352
rect 455418 597408 455474 597417
rect 459560 597382 459612 597388
rect 465078 597408 465134 597417
rect 455418 597343 455474 597352
rect 465078 597343 465134 597352
rect 440240 597314 440292 597320
rect 455432 597310 455460 597343
rect 455420 597304 455472 597310
rect 433338 597272 433394 597281
rect 433338 597207 433394 597216
rect 449898 597272 449954 597281
rect 455420 597246 455472 597252
rect 449898 597207 449900 597216
rect 433352 597174 433380 597207
rect 449952 597207 449954 597216
rect 449900 597178 449952 597184
rect 433340 597168 433392 597174
rect 433340 597110 433392 597116
rect 434718 597136 434774 597145
rect 434718 597071 434720 597080
rect 434772 597071 434774 597080
rect 434720 597042 434772 597048
rect 429200 596896 429252 596902
rect 429200 596838 429252 596844
rect 431958 596864 432014 596873
rect 431958 596799 431960 596808
rect 432012 596799 432014 596808
rect 431960 596770 432012 596776
rect 465092 596766 465120 597343
rect 470598 597000 470654 597009
rect 470598 596935 470600 596944
rect 470652 596935 470654 596944
rect 470600 596906 470652 596912
rect 465080 596760 465132 596766
rect 465080 596702 465132 596708
rect 422574 596456 422630 596465
rect 422574 596391 422630 596400
rect 422588 596358 422616 596391
rect 422576 596352 422628 596358
rect 422576 596294 422628 596300
rect 423678 596320 423734 596329
rect 423678 596255 423680 596264
rect 423732 596255 423734 596264
rect 425058 596320 425114 596329
rect 425058 596255 425114 596264
rect 423680 596226 423732 596232
rect 425072 596222 425100 596255
rect 425060 596216 425112 596222
rect 425060 596158 425112 596164
rect 501604 563100 501656 563106
rect 501604 563042 501656 563048
rect 444380 488776 444432 488782
rect 444380 488718 444432 488724
rect 434720 488708 434772 488714
rect 434720 488650 434772 488656
rect 423680 488504 423732 488510
rect 422574 488472 422630 488481
rect 422574 488407 422576 488416
rect 422628 488407 422630 488416
rect 423678 488472 423680 488481
rect 434732 488481 434760 488650
rect 440240 488572 440292 488578
rect 440240 488514 440292 488520
rect 440252 488481 440280 488514
rect 444392 488481 444420 488718
rect 449900 488640 449952 488646
rect 449900 488582 449952 488588
rect 449912 488481 449940 488582
rect 423732 488472 423734 488481
rect 423678 488407 423734 488416
rect 434718 488472 434774 488481
rect 434718 488407 434774 488416
rect 440238 488472 440294 488481
rect 440238 488407 440294 488416
rect 444378 488472 444434 488481
rect 444378 488407 444434 488416
rect 449898 488472 449954 488481
rect 449898 488407 449954 488416
rect 422576 488378 422628 488384
rect 430578 488336 430634 488345
rect 430578 488271 430634 488280
rect 465078 488336 465134 488345
rect 465078 488271 465134 488280
rect 427818 488200 427874 488209
rect 427818 488135 427820 488144
rect 427872 488135 427874 488144
rect 429198 488200 429254 488209
rect 429198 488135 429254 488144
rect 427820 488106 427872 488112
rect 426438 487792 426494 487801
rect 426438 487727 426440 487736
rect 426492 487727 426494 487736
rect 426440 487698 426492 487704
rect 429212 487626 429240 488135
rect 430592 487694 430620 488271
rect 434718 488200 434774 488209
rect 434718 488135 434774 488144
rect 434732 488102 434760 488135
rect 434720 488096 434772 488102
rect 434720 488038 434772 488044
rect 455418 488064 455474 488073
rect 455418 487999 455474 488008
rect 455432 487966 455460 487999
rect 455420 487960 455472 487966
rect 455420 487902 455472 487908
rect 459558 487928 459614 487937
rect 465092 487898 465120 488271
rect 470598 488064 470654 488073
rect 470598 487999 470600 488008
rect 470652 487999 470654 488008
rect 470600 487970 470652 487976
rect 459558 487863 459614 487872
rect 465080 487892 465132 487898
rect 459572 487830 459600 487863
rect 465080 487834 465132 487840
rect 459560 487824 459612 487830
rect 459560 487766 459612 487772
rect 430580 487688 430632 487694
rect 430580 487630 430632 487636
rect 432050 487656 432106 487665
rect 429200 487620 429252 487626
rect 432050 487591 432106 487600
rect 429200 487562 429252 487568
rect 432064 487558 432092 487591
rect 432052 487552 432104 487558
rect 432052 487494 432104 487500
rect 433338 487384 433394 487393
rect 433338 487319 433394 487328
rect 433352 487286 433380 487319
rect 433340 487280 433392 487286
rect 433340 487222 433392 487228
rect 434718 487248 434774 487257
rect 434718 487183 434720 487192
rect 434772 487183 434774 487192
rect 434720 487154 434772 487160
rect 409144 464500 409196 464506
rect 409144 464442 409196 464448
rect 408040 463140 408092 463146
rect 408040 463082 408092 463088
rect 402244 463072 402296 463078
rect 402244 463014 402296 463020
rect 393964 461848 394016 461854
rect 393964 461790 394016 461796
rect 371516 458924 371568 458930
rect 371516 458866 371568 458872
rect 309048 458856 309100 458862
rect 309048 458798 309100 458804
rect 298836 458788 298888 458794
rect 298836 458730 298888 458736
rect 298744 453484 298796 453490
rect 298744 453426 298796 453432
rect 297548 453348 297600 453354
rect 297548 453290 297600 453296
rect 298006 452432 298062 452441
rect 298006 452367 298062 452376
rect 298020 451314 298048 452367
rect 298008 451308 298060 451314
rect 298008 451250 298060 451256
rect 298848 449206 298876 458730
rect 298928 458652 298980 458658
rect 298928 458594 298980 458600
rect 298940 449274 298968 458594
rect 299572 458584 299624 458590
rect 299572 458526 299624 458532
rect 299020 458380 299072 458386
rect 299020 458322 299072 458328
rect 299032 450566 299060 458322
rect 299584 454714 299612 458526
rect 309060 455940 309088 458798
rect 329656 458788 329708 458794
rect 329656 458730 329708 458736
rect 321284 458516 321336 458522
rect 321284 458458 321336 458464
rect 312912 457292 312964 457298
rect 312912 457234 312964 457240
rect 312924 455940 312952 457234
rect 317420 456272 317472 456278
rect 317420 456214 317472 456220
rect 317432 455940 317460 456214
rect 321296 455940 321324 458458
rect 325792 457224 325844 457230
rect 325792 457166 325844 457172
rect 325804 455940 325832 457166
rect 329668 455940 329696 458730
rect 346400 458720 346452 458726
rect 346400 458662 346452 458668
rect 338028 457156 338080 457162
rect 338028 457098 338080 457104
rect 334164 457020 334216 457026
rect 334164 456962 334216 456968
rect 334176 455940 334204 456962
rect 338040 455940 338068 457098
rect 342536 457088 342588 457094
rect 342536 457030 342588 457036
rect 342548 455940 342576 457030
rect 346412 455940 346440 458662
rect 354772 458652 354824 458658
rect 354772 458594 354824 458600
rect 350908 456952 350960 456958
rect 350908 456894 350960 456900
rect 350920 455940 350948 456894
rect 354784 455940 354812 458594
rect 359280 458584 359332 458590
rect 359280 458526 359332 458532
rect 359292 455940 359320 458526
rect 363144 458448 363196 458454
rect 363144 458390 363196 458396
rect 363156 455940 363184 458390
rect 367652 458380 367704 458386
rect 367652 458322 367704 458328
rect 367664 455940 367692 458322
rect 371528 455940 371556 458866
rect 379888 458312 379940 458318
rect 379888 458254 379940 458260
rect 376024 456884 376076 456890
rect 376024 456826 376076 456832
rect 376036 455940 376064 456826
rect 379900 455940 379928 458254
rect 501616 457502 501644 563042
rect 502996 460358 503024 670686
rect 503076 643136 503128 643142
rect 503076 643078 503128 643084
rect 503088 464438 503116 643078
rect 503168 616888 503220 616894
rect 503168 616830 503220 616836
rect 503076 464432 503128 464438
rect 503076 464374 503128 464380
rect 502984 460352 503036 460358
rect 502984 460294 503036 460300
rect 503180 460290 503208 616830
rect 505756 461718 505784 700266
rect 523684 630692 523736 630698
rect 523684 630634 523736 630640
rect 515404 536852 515456 536858
rect 515404 536794 515456 536800
rect 515416 464370 515444 536794
rect 519544 524476 519596 524482
rect 519544 524418 519596 524424
rect 515404 464364 515456 464370
rect 515404 464306 515456 464312
rect 505744 461712 505796 461718
rect 505744 461654 505796 461660
rect 503168 460284 503220 460290
rect 503168 460226 503220 460232
rect 519556 460222 519584 524418
rect 523696 468586 523724 630634
rect 523684 468580 523736 468586
rect 523684 468522 523736 468528
rect 527192 465730 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 533344 683188 533396 683194
rect 533344 683130 533396 683136
rect 533356 468518 533384 683130
rect 533344 468512 533396 468518
rect 533344 468454 533396 468460
rect 527180 465724 527232 465730
rect 527180 465666 527232 465672
rect 542372 461650 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 549904 510672 549956 510678
rect 549904 510614 549956 510620
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 549916 463010 549944 510614
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580276 467158 580304 577623
rect 580264 467152 580316 467158
rect 580264 467094 580316 467100
rect 549904 463004 549956 463010
rect 549904 462946 549956 462952
rect 542360 461644 542412 461650
rect 542360 461586 542412 461592
rect 519544 460216 519596 460222
rect 519544 460158 519596 460164
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 501604 457496 501656 457502
rect 501604 457438 501656 457444
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 385316 456204 385368 456210
rect 385316 456146 385368 456152
rect 384120 456136 384172 456142
rect 384120 456078 384172 456084
rect 384028 456000 384080 456006
rect 384028 455942 384080 455948
rect 299664 455660 299716 455666
rect 299664 455602 299716 455608
rect 299572 454708 299624 454714
rect 299572 454650 299624 454656
rect 299676 451274 299704 455602
rect 299768 455518 300702 455546
rect 304184 455518 304566 455546
rect 383580 455530 383778 455546
rect 383568 455524 383778 455530
rect 299768 451926 299796 455518
rect 304184 455394 304212 455518
rect 383620 455518 383778 455524
rect 383568 455466 383620 455472
rect 299848 455388 299900 455394
rect 299848 455330 299900 455336
rect 304172 455388 304224 455394
rect 304172 455330 304224 455336
rect 299860 454782 299888 455330
rect 299848 454776 299900 454782
rect 299848 454718 299900 454724
rect 383934 454064 383990 454073
rect 383856 454022 383934 454050
rect 299756 451920 299808 451926
rect 299756 451862 299808 451868
rect 299676 451246 299888 451274
rect 299020 450560 299072 450566
rect 299020 450502 299072 450508
rect 298928 449268 298980 449274
rect 298928 449210 298980 449216
rect 298836 449200 298888 449206
rect 298836 449142 298888 449148
rect 297364 448520 297416 448526
rect 297364 448462 297416 448468
rect 297362 448352 297418 448361
rect 297362 448287 297418 448296
rect 295984 447840 296036 447846
rect 295984 447782 296036 447788
rect 297376 447166 297404 448287
rect 297364 447160 297416 447166
rect 297364 447102 297416 447108
rect 299204 446684 299256 446690
rect 299204 446626 299256 446632
rect 281724 446616 281776 446622
rect 281724 446558 281776 446564
rect 298926 446584 298982 446593
rect 281632 446548 281684 446554
rect 298926 446519 298982 446528
rect 281632 446490 281684 446496
rect 298652 446072 298704 446078
rect 296074 446040 296130 446049
rect 298652 446014 298704 446020
rect 296074 445975 296130 445984
rect 268292 444984 268344 444990
rect 268292 444926 268344 444932
rect 272522 444952 272578 444961
rect 267372 444916 267424 444922
rect 267372 444858 267424 444864
rect 267280 444508 267332 444514
rect 267280 444450 267332 444456
rect 267188 443352 267240 443358
rect 267188 443294 267240 443300
rect 267200 404326 267228 443294
rect 267292 422278 267320 444450
rect 267384 426426 267412 444858
rect 268304 437474 268332 444926
rect 272522 444887 272578 444896
rect 268476 443420 268528 443426
rect 268476 443362 268528 443368
rect 268384 443012 268436 443018
rect 268384 442954 268436 442960
rect 268396 440230 268424 442954
rect 268384 440224 268436 440230
rect 268384 440166 268436 440172
rect 268304 437446 268424 437474
rect 267372 426420 267424 426426
rect 267372 426362 267424 426368
rect 267280 422272 267332 422278
rect 267280 422214 267332 422220
rect 267188 404320 267240 404326
rect 267188 404262 267240 404268
rect 267096 398744 267148 398750
rect 267096 398686 267148 398692
rect 268396 398682 268424 437446
rect 268488 408474 268516 443362
rect 268476 408468 268528 408474
rect 268476 408410 268528 408416
rect 268384 398676 268436 398682
rect 268384 398618 268436 398624
rect 269120 354340 269172 354346
rect 269120 354282 269172 354288
rect 267004 126948 267056 126954
rect 267004 126890 267056 126896
rect 269132 16574 269160 354282
rect 272536 167006 272564 444887
rect 295982 443184 296038 443193
rect 295982 443119 296038 443128
rect 274640 399220 274692 399226
rect 274640 399162 274692 399168
rect 273258 395584 273314 395593
rect 273258 395519 273314 395528
rect 272524 167000 272576 167006
rect 272524 166942 272576 166948
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 261484 9036 261536 9042
rect 261484 8978 261536 8984
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 261772 480 261800 3742
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 265348 6724 265400 6730
rect 265348 6666 265400 6672
rect 264152 3868 264204 3874
rect 264152 3810 264204 3816
rect 264164 480 264192 3810
rect 265360 480 265388 6666
rect 266556 480 266584 16546
rect 268844 7880 268896 7886
rect 268844 7822 268896 7828
rect 267740 6656 267792 6662
rect 267740 6598 267792 6604
rect 267752 480 267780 6598
rect 268856 480 268884 7822
rect 270052 480 270080 16546
rect 272430 9072 272486 9081
rect 272430 9007 272486 9016
rect 271236 6588 271288 6594
rect 271236 6530 271288 6536
rect 271248 480 271276 6530
rect 272444 480 272472 9007
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 395519
rect 274652 16574 274680 399162
rect 282184 398404 282236 398410
rect 282184 398346 282236 398352
rect 277400 392828 277452 392834
rect 277400 392770 277452 392776
rect 276020 24540 276072 24546
rect 276020 24482 276072 24488
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 3806 276060 24482
rect 276110 17504 276166 17513
rect 276110 17439 276166 17448
rect 276020 3800 276072 3806
rect 276020 3742 276072 3748
rect 276124 3482 276152 17439
rect 277412 16574 277440 392770
rect 280160 24472 280212 24478
rect 280160 24414 280212 24420
rect 278780 17672 278832 17678
rect 278780 17614 278832 17620
rect 278792 16574 278820 17614
rect 280172 16574 280200 24414
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276756 3800 276808 3806
rect 276756 3742 276808 3748
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3742
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 282196 6322 282224 398346
rect 289818 396536 289874 396545
rect 289818 396471 289874 396480
rect 284300 354272 284352 354278
rect 284300 354214 284352 354220
rect 282920 17604 282972 17610
rect 282920 17546 282972 17552
rect 282932 16574 282960 17546
rect 282932 16546 283144 16574
rect 281908 6316 281960 6322
rect 281908 6258 281960 6264
rect 282184 6316 282236 6322
rect 282184 6258 282236 6264
rect 281920 480 281948 6258
rect 283116 480 283144 16546
rect 284312 480 284340 354214
rect 285680 84924 285732 84930
rect 285680 84866 285732 84872
rect 285692 16574 285720 84866
rect 287060 26036 287112 26042
rect 287060 25978 287112 25984
rect 287072 16574 287100 25978
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 285404 6520 285456 6526
rect 285404 6462 285456 6468
rect 285416 480 285444 6462
rect 286612 480 286640 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288992 7812 289044 7818
rect 288992 7754 289044 7760
rect 289004 480 289032 7754
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 396471
rect 293960 177744 294012 177750
rect 293960 177686 294012 177692
rect 291198 87680 291254 87689
rect 291198 87615 291254 87624
rect 291212 16574 291240 87615
rect 292578 18592 292634 18601
rect 292578 18527 292634 18536
rect 292592 16574 292620 18527
rect 293972 16574 294000 177686
rect 295996 60722 296024 443119
rect 296088 139398 296116 445975
rect 297364 445868 297416 445874
rect 297364 445810 297416 445816
rect 296536 444848 296588 444854
rect 296536 444790 296588 444796
rect 296444 444780 296496 444786
rect 296444 444722 296496 444728
rect 296352 444712 296404 444718
rect 296352 444654 296404 444660
rect 296260 444644 296312 444650
rect 296260 444586 296312 444592
rect 296166 443320 296222 443329
rect 296166 443255 296222 443264
rect 296076 139392 296128 139398
rect 296076 139334 296128 139340
rect 296180 100706 296208 443255
rect 296272 179382 296300 444586
rect 296364 219434 296392 444654
rect 296456 259418 296484 444722
rect 296548 313274 296576 444790
rect 296626 442232 296682 442241
rect 296626 442167 296682 442176
rect 296640 365702 296668 442167
rect 296996 404320 297048 404326
rect 296996 404262 297048 404268
rect 297008 404161 297036 404262
rect 296994 404152 297050 404161
rect 296994 404087 297050 404096
rect 297376 399430 297404 445810
rect 297640 445120 297692 445126
rect 297640 445062 297692 445068
rect 297548 443692 297600 443698
rect 297548 443634 297600 443640
rect 297456 443556 297508 443562
rect 297456 443498 297508 443504
rect 297364 399424 297416 399430
rect 297364 399366 297416 399372
rect 297468 398546 297496 443498
rect 297560 413001 297588 443634
rect 297652 417081 297680 445062
rect 298006 443592 298062 443601
rect 298006 443527 298062 443536
rect 298020 443086 298048 443527
rect 298560 443284 298612 443290
rect 298560 443226 298612 443232
rect 298008 443080 298060 443086
rect 298008 443022 298060 443028
rect 298008 440224 298060 440230
rect 298008 440166 298060 440172
rect 298020 439521 298048 440166
rect 298006 439512 298062 439521
rect 298006 439447 298062 439456
rect 298008 436076 298060 436082
rect 298008 436018 298060 436024
rect 298020 434761 298048 436018
rect 298006 434752 298062 434761
rect 298006 434687 298062 434696
rect 298008 431928 298060 431934
rect 298008 431870 298060 431876
rect 298020 430681 298048 431870
rect 298006 430672 298062 430681
rect 298006 430607 298062 430616
rect 298008 426420 298060 426426
rect 298008 426362 298060 426368
rect 298020 425921 298048 426362
rect 298006 425912 298062 425921
rect 298006 425847 298062 425856
rect 297916 422272 297968 422278
rect 297916 422214 297968 422220
rect 297928 421841 297956 422214
rect 297914 421832 297970 421841
rect 297914 421767 297970 421776
rect 297638 417072 297694 417081
rect 297638 417007 297694 417016
rect 297546 412992 297602 413001
rect 297546 412927 297602 412936
rect 298008 408468 298060 408474
rect 298008 408410 298060 408416
rect 298020 408241 298048 408410
rect 298006 408232 298062 408241
rect 298006 408167 298062 408176
rect 298572 398614 298600 443226
rect 298664 399226 298692 446014
rect 298836 444576 298888 444582
rect 298836 444518 298888 444524
rect 298742 443728 298798 443737
rect 298742 443663 298798 443672
rect 298652 399220 298704 399226
rect 298652 399162 298704 399168
rect 298560 398608 298612 398614
rect 298560 398550 298612 398556
rect 297456 398540 297508 398546
rect 297456 398482 297508 398488
rect 296628 365696 296680 365702
rect 296628 365638 296680 365644
rect 296536 313268 296588 313274
rect 296536 313210 296588 313216
rect 296444 259412 296496 259418
rect 296444 259354 296496 259360
rect 296352 219428 296404 219434
rect 296352 219370 296404 219376
rect 298756 193186 298784 443663
rect 298848 245614 298876 444518
rect 298940 273222 298968 446519
rect 299020 445936 299072 445942
rect 299020 445878 299072 445884
rect 299032 325650 299060 445878
rect 299112 443148 299164 443154
rect 299112 443090 299164 443096
rect 299124 379506 299152 443090
rect 299216 398818 299244 446626
rect 299860 446418 299888 451246
rect 299848 446412 299900 446418
rect 299848 446354 299900 446360
rect 299388 446140 299440 446146
rect 299388 446082 299440 446088
rect 299296 446004 299348 446010
rect 299296 445946 299348 445952
rect 299308 400178 299336 445946
rect 299296 400172 299348 400178
rect 299296 400114 299348 400120
rect 299400 399294 299428 446082
rect 299480 445052 299532 445058
rect 299480 444994 299532 445000
rect 299492 422294 299520 444994
rect 383856 431954 383884 454022
rect 383934 453999 383990 454008
rect 384040 452305 384068 455942
rect 384026 452296 384082 452305
rect 384026 452231 384082 452240
rect 384132 452146 384160 456078
rect 384212 456068 384264 456074
rect 384212 456010 384264 456016
rect 383948 452118 384160 452146
rect 383948 438705 383976 452118
rect 384224 451274 384252 456010
rect 385040 455932 385092 455938
rect 385040 455874 385092 455880
rect 384304 455592 384356 455598
rect 384304 455534 384356 455540
rect 384040 451246 384252 451274
rect 384040 448225 384068 451246
rect 384026 448216 384082 448225
rect 384026 448151 384082 448160
rect 383934 438696 383990 438705
rect 383934 438631 383990 438640
rect 383856 431926 383976 431954
rect 384316 431934 384344 455534
rect 299492 422266 299704 422294
rect 299676 400738 299704 422266
rect 383948 421705 383976 431926
rect 384304 431928 384356 431934
rect 384304 431870 384356 431876
rect 383934 421696 383990 421705
rect 383934 421631 383990 421640
rect 385052 412321 385080 455874
rect 385224 455796 385276 455802
rect 385224 455738 385276 455744
rect 385132 455660 385184 455666
rect 385132 455602 385184 455608
rect 385144 416401 385172 455602
rect 385236 425241 385264 455738
rect 385328 430001 385356 456146
rect 385408 455864 385460 455870
rect 385408 455806 385460 455812
rect 385420 434081 385448 455806
rect 385500 455728 385552 455734
rect 385500 455670 385552 455676
rect 385512 442921 385540 455670
rect 580264 455456 580316 455462
rect 580264 455398 580316 455404
rect 385498 442912 385554 442921
rect 385498 442847 385554 442856
rect 385406 434072 385462 434081
rect 385406 434007 385462 434016
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 385314 429992 385370 430001
rect 385314 429927 385370 429936
rect 385222 425232 385278 425241
rect 385222 425167 385278 425176
rect 580276 418305 580304 455398
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 385130 416392 385186 416401
rect 385130 416327 385186 416336
rect 385038 412312 385094 412321
rect 385038 412247 385094 412256
rect 385038 407552 385094 407561
rect 385038 407487 385094 407496
rect 385052 401266 385080 407487
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 385040 401260 385092 401266
rect 385040 401202 385092 401208
rect 299676 400710 300058 400738
rect 328840 400722 329038 400738
rect 370608 400722 370898 400738
rect 328828 400716 329038 400722
rect 328880 400710 329038 400716
rect 370596 400716 370898 400722
rect 328828 400658 328880 400664
rect 370648 400710 370898 400716
rect 370596 400658 370648 400664
rect 580000 400178 580028 404903
rect 579988 400172 580040 400178
rect 579988 400114 580040 400120
rect 299388 399288 299440 399294
rect 299388 399230 299440 399236
rect 303908 398818 303936 400044
rect 307772 399430 307800 400044
rect 307760 399424 307812 399430
rect 307760 399366 307812 399372
rect 312280 399129 312308 400044
rect 312266 399120 312322 399129
rect 312266 399055 312322 399064
rect 299204 398812 299256 398818
rect 299204 398754 299256 398760
rect 303896 398812 303948 398818
rect 303896 398754 303948 398760
rect 316144 398313 316172 400044
rect 320652 398546 320680 400044
rect 324516 399129 324544 400044
rect 331220 399492 331272 399498
rect 331220 399434 331272 399440
rect 324502 399120 324558 399129
rect 324502 399055 324558 399064
rect 320640 398540 320692 398546
rect 320640 398482 320692 398488
rect 316130 398304 316186 398313
rect 316130 398239 316186 398248
rect 310518 397352 310574 397361
rect 310518 397287 310574 397296
rect 307760 396908 307812 396914
rect 307760 396850 307812 396856
rect 300860 389836 300912 389842
rect 300860 389778 300912 389784
rect 299112 379500 299164 379506
rect 299112 379442 299164 379448
rect 299020 325644 299072 325650
rect 299020 325586 299072 325592
rect 298928 273216 298980 273222
rect 298928 273158 298980 273164
rect 298836 245608 298888 245614
rect 298836 245550 298888 245556
rect 298744 193180 298796 193186
rect 298744 193122 298796 193128
rect 296260 179376 296312 179382
rect 296260 179318 296312 179324
rect 298100 177676 298152 177682
rect 298100 177618 298152 177624
rect 296168 100700 296220 100706
rect 296168 100642 296220 100648
rect 295984 60716 296036 60722
rect 295984 60658 296036 60664
rect 296720 19100 296772 19106
rect 296720 19042 296772 19048
rect 296732 16574 296760 19042
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 291396 480 291424 16546
rect 292578 7848 292634 7857
rect 292578 7783 292634 7792
rect 292592 480 292620 7783
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 296076 3732 296128 3738
rect 296076 3674 296128 3680
rect 296088 480 296116 3674
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 177618
rect 299480 19032 299532 19038
rect 299480 18974 299532 18980
rect 299492 3398 299520 18974
rect 300872 16574 300900 389778
rect 304998 354376 305054 354385
rect 304998 354311 305054 354320
rect 303620 18964 303672 18970
rect 303620 18906 303672 18912
rect 303632 16574 303660 18906
rect 305012 16574 305040 354311
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299662 3768 299718 3777
rect 299662 3703 299718 3712
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 299676 480 299704 3703
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303160 7744 303212 7750
rect 303160 7686 303212 7692
rect 303172 480 303200 7686
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306746 7712 306802 7721
rect 306746 7647 306802 7656
rect 306760 480 306788 7647
rect 307772 3482 307800 396850
rect 307852 394460 307904 394466
rect 307852 394402 307904 394408
rect 307864 3738 307892 394402
rect 310532 16574 310560 397287
rect 324318 397216 324374 397225
rect 324318 397151 324374 397160
rect 318800 394392 318852 394398
rect 318800 394334 318852 394340
rect 313280 391536 313332 391542
rect 313280 391478 313332 391484
rect 311900 25968 311952 25974
rect 311900 25910 311952 25916
rect 311912 16574 311940 25910
rect 313292 16574 313320 391478
rect 316040 355700 316092 355706
rect 316040 355642 316092 355648
rect 314660 18896 314712 18902
rect 314660 18838 314712 18844
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 310242 7576 310298 7585
rect 310242 7511 310298 7520
rect 307852 3732 307904 3738
rect 307852 3674 307904 3680
rect 309048 3732 309100 3738
rect 309048 3674 309100 3680
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 3674
rect 310256 480 310284 7511
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 18838
rect 316052 3482 316080 355642
rect 316132 87780 316184 87786
rect 316132 87722 316184 87728
rect 316144 3738 316172 87722
rect 317420 18828 317472 18834
rect 317420 18770 317472 18776
rect 317432 16574 317460 18770
rect 318812 16574 318840 394334
rect 322940 25900 322992 25906
rect 322940 25842 322992 25848
rect 321560 18760 321612 18766
rect 321560 18702 321612 18708
rect 321572 16574 321600 18702
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 321572 16546 322152 16574
rect 316132 3732 316184 3738
rect 316132 3674 316184 3680
rect 317328 3732 317380 3738
rect 317328 3674 317380 3680
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 3674
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 320916 9444 320968 9450
rect 320916 9386 320968 9392
rect 320928 480 320956 9386
rect 322124 480 322152 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 25842
rect 324332 3398 324360 397151
rect 328458 397080 328514 397089
rect 328458 397015 328514 397024
rect 325698 393952 325754 393961
rect 325698 393887 325754 393896
rect 324412 355632 324464 355638
rect 324412 355574 324464 355580
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 355574
rect 325712 16574 325740 393887
rect 328472 16574 328500 397015
rect 329840 394324 329892 394330
rect 329840 394266 329892 394272
rect 329852 16574 329880 394266
rect 325712 16546 326384 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 327998 8936 328054 8945
rect 327998 8871 328054 8880
rect 328012 480 328040 8871
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 399434
rect 332888 398449 332916 400044
rect 333980 399356 334032 399362
rect 333980 399298 334032 399304
rect 332874 398440 332930 398449
rect 332874 398375 332930 398384
rect 332600 25832 332652 25838
rect 332600 25774 332652 25780
rect 332612 3398 332640 25774
rect 332692 18692 332744 18698
rect 332692 18634 332744 18640
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 18634
rect 333992 16574 334020 399298
rect 337396 399158 337424 400044
rect 341260 399294 341288 400044
rect 341248 399288 341300 399294
rect 341248 399230 341300 399236
rect 337384 399152 337436 399158
rect 337384 399094 337436 399100
rect 345768 399090 345796 400044
rect 345756 399084 345808 399090
rect 345756 399026 345808 399032
rect 349632 398614 349660 400044
rect 354140 398682 354168 400044
rect 354128 398676 354180 398682
rect 354128 398618 354180 398624
rect 349620 398608 349672 398614
rect 358004 398585 358032 400044
rect 362512 398721 362540 400044
rect 366376 399226 366404 400044
rect 366364 399220 366416 399226
rect 366364 399162 366416 399168
rect 374748 398750 374776 400044
rect 379256 398857 379284 400044
rect 379242 398848 379298 398857
rect 379242 398783 379298 398792
rect 374736 398744 374788 398750
rect 362498 398712 362554 398721
rect 374736 398686 374788 398692
rect 362498 398647 362554 398656
rect 349620 398550 349672 398556
rect 357990 398576 358046 398585
rect 357990 398511 358046 398520
rect 383120 398342 383148 400044
rect 580262 399528 580318 399537
rect 580262 399463 580318 399472
rect 383660 399016 383712 399022
rect 383660 398958 383712 398964
rect 383108 398336 383160 398342
rect 383108 398278 383160 398284
rect 364338 396944 364394 396953
rect 364338 396879 364394 396888
rect 339500 396840 339552 396846
rect 339500 396782 339552 396788
rect 336740 23180 336792 23186
rect 336740 23122 336792 23128
rect 335360 18624 335412 18630
rect 335360 18566 335412 18572
rect 335372 16574 335400 18566
rect 336752 16574 336780 23122
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338672 9376 338724 9382
rect 338672 9318 338724 9324
rect 338684 480 338712 9318
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 396782
rect 340880 394256 340932 394262
rect 340880 394198 340932 394204
rect 340892 16574 340920 394198
rect 347780 394188 347832 394194
rect 347780 394130 347832 394136
rect 345018 355600 345074 355609
rect 345018 355535 345074 355544
rect 342260 351280 342312 351286
rect 342260 351222 342312 351228
rect 342272 16574 342300 351222
rect 343638 25528 343694 25537
rect 343638 25463 343694 25472
rect 343652 16574 343680 25463
rect 345032 16574 345060 355535
rect 346398 353016 346454 353025
rect 346398 352951 346454 352960
rect 346412 16574 346440 352951
rect 347792 16574 347820 394130
rect 349160 392760 349212 392766
rect 349160 392702 349212 392708
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 340984 480 341012 16546
rect 342168 9308 342220 9314
rect 342168 9250 342220 9256
rect 342180 480 342208 9250
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 392702
rect 350540 356720 350592 356726
rect 350540 356662 350592 356668
rect 349252 20256 349304 20262
rect 349252 20198 349304 20204
rect 349264 3398 349292 20198
rect 350552 16574 350580 356662
rect 357440 355564 357492 355570
rect 357440 355506 357492 355512
rect 353300 20188 353352 20194
rect 353300 20130 353352 20136
rect 353312 16574 353340 20130
rect 350552 16546 351224 16574
rect 353312 16546 353616 16574
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352840 9240 352892 9246
rect 352840 9182 352892 9188
rect 352852 480 352880 9182
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 356336 9172 356388 9178
rect 356336 9114 356388 9120
rect 355232 5160 355284 5166
rect 355232 5102 355284 5108
rect 355244 480 355272 5102
rect 356348 480 356376 9114
rect 357452 3398 357480 355506
rect 360198 355464 360254 355473
rect 360198 355399 360254 355408
rect 357532 354204 357584 354210
rect 357532 354146 357584 354152
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 354146
rect 360212 16574 360240 355399
rect 364352 16574 364380 396879
rect 372620 395752 372672 395758
rect 372620 395694 372672 395700
rect 365720 394120 365772 394126
rect 365720 394062 365772 394068
rect 360212 16546 361160 16574
rect 364352 16546 364656 16574
rect 359924 9104 359976 9110
rect 359924 9046 359976 9052
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 359936 480 359964 9046
rect 361132 480 361160 16546
rect 363510 10568 363566 10577
rect 363510 10503 363566 10512
rect 362314 5128 362370 5137
rect 362314 5063 362370 5072
rect 362328 480 362356 5063
rect 363524 480 363552 10503
rect 364628 480 364656 16546
rect 365732 3210 365760 394062
rect 368480 394052 368532 394058
rect 368480 393994 368532 394000
rect 367100 355496 367152 355502
rect 367100 355438 367152 355444
rect 367112 16574 367140 355438
rect 368492 16574 368520 393994
rect 371240 355428 371292 355434
rect 371240 355370 371292 355376
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 365812 10668 365864 10674
rect 365812 10610 365864 10616
rect 365824 3398 365852 10610
rect 365812 3392 365864 3398
rect 365812 3334 365864 3340
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 365732 3182 365852 3210
rect 365824 480 365852 3182
rect 367020 480 367048 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370136 10600 370188 10606
rect 370136 10542 370188 10548
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 10542
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 355370
rect 372632 16574 372660 395694
rect 379520 393984 379572 393990
rect 379520 393926 379572 393932
rect 375380 25764 375432 25770
rect 375380 25706 375432 25712
rect 374000 20120 374052 20126
rect 374000 20062 374052 20068
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3398 374040 20062
rect 375392 16574 375420 25706
rect 378138 20224 378194 20233
rect 378138 20159 378194 20168
rect 378152 16574 378180 20159
rect 375392 16546 376064 16574
rect 378152 16546 378456 16574
rect 374092 10532 374144 10538
rect 374092 10474 374144 10480
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 10474
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377678 10432 377734 10441
rect 377678 10367 377734 10376
rect 377692 480 377720 10367
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 393926
rect 382280 177608 382332 177614
rect 382280 177550 382332 177556
rect 381174 10296 381230 10305
rect 381174 10231 381230 10240
rect 381188 480 381216 10231
rect 382292 3398 382320 177550
rect 382370 20088 382426 20097
rect 382370 20023 382426 20032
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 20023
rect 383672 16574 383700 398958
rect 400220 398948 400272 398954
rect 400220 398890 400272 398896
rect 396080 396772 396132 396778
rect 396080 396714 396132 396720
rect 385040 391468 385092 391474
rect 385040 391410 385092 391416
rect 385052 16574 385080 391410
rect 393320 355360 393372 355366
rect 393320 355302 393372 355308
rect 386420 228404 386472 228410
rect 386420 228346 386472 228352
rect 386432 16574 386460 228346
rect 390560 177540 390612 177546
rect 390560 177482 390612 177488
rect 389180 20052 389232 20058
rect 389180 19994 389232 20000
rect 389192 16574 389220 19994
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387800 10464 387852 10470
rect 387800 10406 387852 10412
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 10406
rect 389468 480 389496 16546
rect 390572 3210 390600 177482
rect 391940 19984 391992 19990
rect 391940 19926 391992 19932
rect 391952 16574 391980 19926
rect 393332 16574 393360 355302
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 390652 10396 390704 10402
rect 390652 10338 390704 10344
rect 390664 3398 390692 10338
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395344 12096 395396 12102
rect 395344 12038 395396 12044
rect 395356 480 395384 12038
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 396714
rect 397460 354136 397512 354142
rect 397460 354078 397512 354084
rect 397472 16574 397500 354078
rect 398838 351248 398894 351257
rect 398838 351183 398894 351192
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3398 398880 351183
rect 400232 16574 400260 398890
rect 455420 398880 455472 398886
rect 455420 398822 455472 398828
rect 416778 396808 416834 396817
rect 416778 396743 416834 396752
rect 414018 352880 414074 352889
rect 414018 352815 414074 352824
rect 407120 87712 407172 87718
rect 407120 87654 407172 87660
rect 402980 83496 403032 83502
rect 402980 83438 403032 83444
rect 402992 16574 403020 83438
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 398930 11928 398986 11937
rect 398930 11863 398986 11872
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 11863
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 12028 402572 12034
rect 402520 11970 402572 11976
rect 402532 480 402560 11970
rect 403636 480 403664 16546
rect 406016 11960 406068 11966
rect 406016 11902 406068 11908
rect 404820 6452 404872 6458
rect 404820 6394 404872 6400
rect 404832 480 404860 6394
rect 406028 480 406056 11902
rect 407132 3210 407160 87654
rect 407212 26988 407264 26994
rect 407212 26930 407264 26936
rect 407224 3398 407252 26930
rect 409880 21888 409932 21894
rect 409880 21830 409932 21836
rect 409892 16574 409920 21830
rect 414032 16574 414060 352815
rect 415400 26920 415452 26926
rect 415400 26862 415452 26868
rect 409892 16546 410840 16574
rect 414032 16546 414336 16574
rect 409144 11892 409196 11898
rect 409144 11834 409196 11840
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 11834
rect 410812 480 410840 16546
rect 412638 11792 412694 11801
rect 412638 11727 412694 11736
rect 411904 6384 411956 6390
rect 411904 6326 411956 6332
rect 411916 480 411944 6326
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 11727
rect 414308 480 414336 16546
rect 415412 3210 415440 26862
rect 416792 16574 416820 396743
rect 445760 392692 445812 392698
rect 445760 392634 445812 392640
rect 419540 391400 419592 391406
rect 419540 391342 419592 391348
rect 419552 16574 419580 391342
rect 437480 391332 437532 391338
rect 437480 391274 437532 391280
rect 431958 354240 432014 354249
rect 431958 354175 432014 354184
rect 425060 25696 425112 25702
rect 425060 25638 425112 25644
rect 420920 21820 420972 21826
rect 420920 21762 420972 21768
rect 416792 16546 417464 16574
rect 419552 16546 420224 16574
rect 415490 11656 415546 11665
rect 415490 11591 415546 11600
rect 415504 3398 415532 11591
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 3182 415532 3210
rect 415504 480 415532 3182
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418528 16312 418580 16318
rect 418528 16254 418580 16260
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16254
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 21762
rect 423680 21752 423732 21758
rect 423680 21694 423732 21700
rect 422576 7676 422628 7682
rect 422576 7618 422628 7624
rect 422588 480 422616 7618
rect 423692 1698 423720 21694
rect 425072 16574 425100 25638
rect 427820 21684 427872 21690
rect 427820 21626 427872 21632
rect 427832 16574 427860 21626
rect 425072 16546 425744 16574
rect 427832 16546 428504 16574
rect 423772 11824 423824 11830
rect 423772 11766 423824 11772
rect 423680 1692 423732 1698
rect 423680 1634 423732 1640
rect 423784 480 423812 11766
rect 424968 1692 425020 1698
rect 424968 1634 425020 1640
rect 424980 480 425008 1634
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426808 11756 426860 11762
rect 426808 11698 426860 11704
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 11698
rect 428476 480 428504 16546
rect 430856 13524 430908 13530
rect 430856 13466 430908 13472
rect 429660 7608 429712 7614
rect 429660 7550 429712 7556
rect 429672 480 429700 7550
rect 430868 480 430896 13466
rect 431972 1170 432000 354175
rect 436100 352708 436152 352714
rect 436100 352650 436152 352656
rect 432050 87544 432106 87553
rect 432050 87479 432106 87488
rect 432064 3398 432092 87479
rect 434718 21312 434774 21321
rect 434718 21247 434774 21256
rect 434732 16574 434760 21247
rect 436112 16574 436140 352650
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433982 13152 434038 13161
rect 433982 13087 434038 13096
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 13087
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 391274
rect 443000 35216 443052 35222
rect 443000 35158 443052 35164
rect 440240 25628 440292 25634
rect 440240 25570 440292 25576
rect 438860 21616 438912 21622
rect 438860 21558 438912 21564
rect 438872 16574 438900 21558
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 25570
rect 441620 21548 441672 21554
rect 441620 21490 441672 21496
rect 441632 16574 441660 21490
rect 443012 16574 443040 35158
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 440332 13456 440384 13462
rect 440332 13398 440384 13404
rect 440344 3398 440372 13398
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445024 13388 445076 13394
rect 445024 13330 445076 13336
rect 445036 480 445064 13330
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 392634
rect 452658 354104 452714 354113
rect 452658 354039 452714 354048
rect 449900 302932 449952 302938
rect 449900 302874 449952 302880
rect 448520 87644 448572 87650
rect 448520 87586 448572 87592
rect 447140 25560 447192 25566
rect 447140 25502 447192 25508
rect 447152 16574 447180 25502
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 1698 448560 87586
rect 449912 16574 449940 302874
rect 452672 16574 452700 354039
rect 454040 49020 454092 49026
rect 454040 48962 454092 48968
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 448612 13320 448664 13326
rect 448612 13262 448664 13268
rect 448520 1692 448572 1698
rect 448520 1634 448572 1640
rect 448624 480 448652 13262
rect 449808 1692 449860 1698
rect 449808 1634 449860 1640
rect 449820 480 449848 1634
rect 450924 480 450952 16546
rect 451646 13016 451702 13025
rect 451646 12951 451702 12960
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 12951
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 48962
rect 455432 16574 455460 398822
rect 543740 398200 543792 398206
rect 489918 398168 489974 398177
rect 543740 398142 543792 398148
rect 489918 398103 489974 398112
rect 480260 392624 480312 392630
rect 480260 392566 480312 392572
rect 460940 336048 460992 336054
rect 460940 335990 460992 335996
rect 456892 21480 456944 21486
rect 456892 21422 456944 21428
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456904 480 456932 21422
rect 459560 21412 459612 21418
rect 459560 21354 459612 21360
rect 459572 16574 459600 21354
rect 460952 16574 460980 335990
rect 467840 182844 467892 182850
rect 467840 182786 467892 182792
rect 465078 26888 465134 26897
rect 465078 26823 465134 26832
rect 463700 23112 463752 23118
rect 463700 23054 463752 23060
rect 463712 16574 463740 23054
rect 465092 16574 465120 26823
rect 466458 22808 466514 22817
rect 466458 22743 466514 22752
rect 466472 16574 466500 22743
rect 467852 16574 467880 182786
rect 478880 177472 478932 177478
rect 478880 177414 478932 177420
rect 477500 82136 477552 82142
rect 477500 82078 477552 82084
rect 473360 23044 473412 23050
rect 473360 22986 473412 22992
rect 470598 19952 470654 19961
rect 470598 19887 470654 19896
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 465092 16546 465212 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 459192 13252 459244 13258
rect 459192 13194 459244 13200
rect 458088 3664 458140 3670
rect 458088 3606 458140 3612
rect 458100 480 458128 3606
rect 459204 480 459232 13194
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 462320 13184 462372 13190
rect 462320 13126 462372 13132
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 13126
rect 463988 480 464016 16546
rect 465184 480 465212 16546
rect 465816 13116 465868 13122
rect 465816 13058 465868 13064
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 13058
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469862 14784 469918 14793
rect 469862 14719 469918 14728
rect 469876 480 469904 14719
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 19887
rect 473372 3602 473400 22986
rect 477512 16574 477540 82078
rect 477512 16546 478184 16574
rect 473452 14816 473504 14822
rect 473452 14758 473504 14764
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 473360 3596 473412 3602
rect 473360 3538 473412 3544
rect 472268 480 472296 3538
rect 473464 480 473492 14758
rect 476488 14748 476540 14754
rect 476488 14690 476540 14696
rect 475752 9036 475804 9042
rect 475752 8978 475804 8984
rect 474188 3596 474240 3602
rect 474188 3538 474240 3544
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3538
rect 475764 480 475792 8978
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 14690
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 177414
rect 480272 16574 480300 392566
rect 485778 352744 485834 352753
rect 485778 352679 485834 352688
rect 481640 86352 481692 86358
rect 481640 86294 481692 86300
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 3534 481680 86294
rect 485792 16574 485820 352679
rect 485792 16546 486464 16574
rect 481732 14680 481784 14686
rect 481732 14622 481784 14628
rect 484766 14648 484822 14657
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 14622
rect 484766 14583 484822 14592
rect 484032 3596 484084 3602
rect 484032 3538 484084 3544
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 3538
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 14583
rect 486436 480 486464 16546
rect 488814 14512 488870 14521
rect 488814 14447 488870 14456
rect 487618 3632 487674 3641
rect 487618 3567 487674 3576
rect 487632 480 487660 3567
rect 488828 480 488856 14447
rect 489932 3534 489960 398103
rect 507858 398032 507914 398041
rect 507858 397967 507914 397976
rect 499580 395684 499632 395690
rect 499580 395626 499632 395632
rect 492680 391264 492732 391270
rect 492680 391206 492732 391212
rect 490012 22976 490064 22982
rect 490012 22918 490064 22924
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 22918
rect 492692 16574 492720 391206
rect 494060 28348 494112 28354
rect 494060 28290 494112 28296
rect 494072 16574 494100 28290
rect 498200 28280 498252 28286
rect 498200 28222 498252 28228
rect 496820 22908 496872 22914
rect 496820 22850 496872 22856
rect 496832 16574 496860 22850
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 492312 14612 492364 14618
rect 492312 14554 492364 14560
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 14554
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 495440 14544 495492 14550
rect 495440 14486 495492 14492
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 14486
rect 497108 480 497136 16546
rect 498212 480 498240 28222
rect 499592 16574 499620 395626
rect 506478 355328 506534 355337
rect 506478 355263 506534 355272
rect 502340 89004 502392 89010
rect 502340 88946 502392 88952
rect 502352 16574 502380 88946
rect 503718 22672 503774 22681
rect 503718 22607 503774 22616
rect 499592 16546 500632 16574
rect 502352 16546 503024 16574
rect 498936 16244 498988 16250
rect 498936 16186 498988 16192
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16186
rect 500604 480 500632 16546
rect 501788 5092 501840 5098
rect 501788 5034 501840 5040
rect 501800 480 501828 5034
rect 502996 480 503024 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 22607
rect 505374 4992 505430 5001
rect 505374 4927 505430 4936
rect 505388 480 505416 4927
rect 506492 480 506520 355263
rect 506572 22840 506624 22846
rect 506572 22782 506624 22788
rect 506584 16574 506612 22782
rect 507872 16574 507900 397967
rect 525800 397656 525852 397662
rect 525800 397598 525852 397604
rect 514760 395616 514812 395622
rect 514760 395558 514812 395564
rect 512000 352640 512052 352646
rect 512000 352582 512052 352588
rect 510620 22772 510672 22778
rect 510620 22714 510672 22720
rect 510632 16574 510660 22714
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 509608 16176 509660 16182
rect 509608 16118 509660 16124
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16118
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 352582
rect 513380 16108 513432 16114
rect 513380 16050 513432 16056
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 16050
rect 514772 480 514800 395558
rect 521658 395448 521714 395457
rect 521658 395383 521714 395392
rect 518900 177404 518952 177410
rect 518900 177346 518952 177352
rect 514852 86284 514904 86290
rect 514852 86226 514904 86232
rect 514864 16574 514892 86226
rect 517520 24404 517572 24410
rect 517520 24346 517572 24352
rect 517532 16574 517560 24346
rect 518912 16574 518940 177346
rect 514864 16546 515536 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517152 16040 517204 16046
rect 517152 15982 517204 15988
rect 517164 480 517192 15982
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 520278 16008 520334 16017
rect 520278 15943 520334 15952
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 15943
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 395383
rect 524420 352572 524472 352578
rect 524420 352514 524472 352520
rect 524432 16574 524460 352514
rect 525812 16574 525840 397598
rect 528560 395548 528612 395554
rect 528560 395490 528612 395496
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523774 15872 523830 15881
rect 523774 15807 523830 15816
rect 523038 3496 523094 3505
rect 523038 3431 523094 3440
rect 523052 480 523080 3431
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 15807
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 15972 527876 15978
rect 527824 15914 527876 15920
rect 527836 480 527864 15914
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 395490
rect 535460 395480 535512 395486
rect 535460 395422 535512 395428
rect 531320 354068 531372 354074
rect 531320 354010 531372 354016
rect 531332 3534 531360 354010
rect 532700 177336 532752 177342
rect 532700 177278 532752 177284
rect 532712 16574 532740 177278
rect 534080 17536 534132 17542
rect 534080 17478 534132 17484
rect 534092 16574 534120 17478
rect 535472 16574 535500 395422
rect 540978 352608 541034 352617
rect 540978 352543 541034 352552
rect 538218 351112 538274 351121
rect 538218 351047 538274 351056
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 531412 15904 531464 15910
rect 531412 15846 531464 15852
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 530124 3460 530176 3466
rect 530124 3402 530176 3408
rect 530136 480 530164 3402
rect 531424 3346 531452 15846
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 5024 537260 5030
rect 537208 4966 537260 4972
rect 537220 480 537248 4966
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 351047
rect 539598 24304 539654 24313
rect 539598 24239 539654 24248
rect 539612 480 539640 24239
rect 540992 16574 541020 352543
rect 542360 24336 542412 24342
rect 542360 24278 542412 24284
rect 542372 16574 542400 24278
rect 543752 16574 543780 398142
rect 561680 398132 561732 398138
rect 561680 398074 561732 398080
rect 549260 395412 549312 395418
rect 549260 395354 549312 395360
rect 546500 24268 546552 24274
rect 546500 24210 546552 24216
rect 545120 17468 545172 17474
rect 545120 17410 545172 17416
rect 545132 16574 545160 17410
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540794 4856 540850 4865
rect 540794 4791 540850 4800
rect 540808 480 540836 4791
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 24210
rect 547880 17400 547932 17406
rect 547880 17342 547932 17348
rect 547892 16574 547920 17342
rect 549272 16574 549300 395354
rect 556158 395312 556214 395321
rect 556158 395247 556214 395256
rect 554780 351212 554832 351218
rect 554780 351154 554832 351160
rect 553400 24200 553452 24206
rect 553400 24142 553452 24148
rect 552020 17332 552072 17338
rect 552020 17274 552072 17280
rect 552032 16574 552060 17274
rect 553412 16574 553440 24142
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 547880 4956 547932 4962
rect 547880 4898 547932 4904
rect 547892 480 547920 4898
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 551468 4888 551520 4894
rect 551468 4830 551520 4836
rect 551480 480 551508 4830
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 351154
rect 556172 3534 556200 395247
rect 560300 354000 560352 354006
rect 557538 353968 557594 353977
rect 560300 353942 560352 353948
rect 557538 353903 557594 353912
rect 556250 17368 556306 17377
rect 556250 17303 556306 17312
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 17303
rect 557552 16574 557580 353903
rect 558918 17232 558974 17241
rect 558918 17167 558974 17176
rect 558932 16574 558960 17167
rect 560312 16574 560340 353942
rect 561692 16574 561720 398074
rect 564440 397588 564492 397594
rect 564440 397530 564492 397536
rect 563060 84856 563112 84862
rect 563060 84798 563112 84804
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 84798
rect 564452 3534 564480 397530
rect 576858 396672 576914 396681
rect 576858 396607 576914 396616
rect 571340 395344 571392 395350
rect 571340 395286 571392 395292
rect 564532 24132 564584 24138
rect 564532 24074 564584 24080
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 24074
rect 567200 17264 567252 17270
rect 567200 17206 567252 17212
rect 567212 16574 567240 17206
rect 567212 16546 567608 16574
rect 566832 8968 566884 8974
rect 566832 8910 566884 8916
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 8910
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 570328 14476 570380 14482
rect 570328 14418 570380 14424
rect 569132 6248 569184 6254
rect 569132 6190 569184 6196
rect 569144 480 569172 6190
rect 570340 480 570368 14418
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 395286
rect 572720 347064 572772 347070
rect 572720 347006 572772 347012
rect 572732 16574 572760 347006
rect 574098 24168 574154 24177
rect 574098 24103 574154 24112
rect 574112 16574 574140 24103
rect 576872 16574 576900 396607
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580276 152697 580304 399463
rect 582380 397520 582432 397526
rect 582380 397462 582432 397468
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580264 58676 580316 58682
rect 580264 58618 580316 58624
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 572720 6180 572772 6186
rect 572720 6122 572772 6128
rect 572732 480 572760 6122
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576306 6216 576362 6225
rect 576306 6151 576362 6160
rect 576320 480 576348 6151
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 580276 6633 580304 58618
rect 582392 16574 582420 397462
rect 582392 16546 583432 16574
rect 581736 10328 581788 10334
rect 581736 10270 581788 10276
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 6316 581052 6322
rect 581000 6258 581052 6264
rect 578608 4820 578660 4826
rect 578608 4762 578660 4768
rect 578620 480 578648 4762
rect 579802 3360 579858 3369
rect 579802 3295 579858 3304
rect 579816 480 579844 3295
rect 581012 480 581040 6258
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 10270
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 2778 658144 2834 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 619112 3478 619168
rect 3146 606056 3202 606112
rect 2778 579964 2834 580000
rect 2778 579944 2780 579964
rect 2780 579944 2832 579964
rect 2832 579944 2834 579964
rect 3330 553832 3386 553888
rect 2778 527856 2834 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3330 501744 3386 501800
rect 3054 475632 3110 475688
rect 3514 566888 3570 566944
rect 3422 462576 3478 462632
rect 2870 449520 2926 449576
rect 78586 636384 78642 636440
rect 78310 635296 78366 635352
rect 78218 633664 78274 633720
rect 77942 632576 77998 632632
rect 77758 629584 77814 629640
rect 77574 523232 77630 523288
rect 77850 608640 77906 608696
rect 77758 520240 77814 520296
rect 77666 498344 77722 498400
rect 78126 630944 78182 631000
rect 78034 627952 78090 628008
rect 78402 610000 78458 610056
rect 78586 607688 78642 607744
rect 103150 597488 103206 597544
rect 111706 597488 111762 597544
rect 115846 597524 115848 597544
rect 115848 597524 115900 597544
rect 115900 597524 115902 597544
rect 115846 597488 115902 597524
rect 121366 597488 121422 597544
rect 126886 597508 126942 597544
rect 126886 597488 126888 597508
rect 126888 597488 126940 597508
rect 126940 597488 126942 597508
rect 92478 597352 92534 597408
rect 94042 597080 94098 597136
rect 103426 597080 103482 597136
rect 106186 597100 106242 597136
rect 106186 597080 106188 597100
rect 106188 597080 106240 597100
rect 106240 597080 106242 597100
rect 78494 526632 78550 526688
rect 78310 526496 78366 526552
rect 78310 523640 78366 523696
rect 77942 523232 77998 523288
rect 78126 520920 78182 520976
rect 78034 517928 78090 517984
rect 77942 498616 77998 498672
rect 78586 499840 78642 499896
rect 100666 596964 100722 597000
rect 100666 596944 100668 596964
rect 100668 596944 100720 596964
rect 100720 596944 100722 596964
rect 131026 597488 131082 597544
rect 136546 597488 136602 597544
rect 140686 597488 140742 597544
rect 104806 596828 104862 596864
rect 104806 596808 104808 596828
rect 104808 596808 104860 596828
rect 104860 596808 104862 596828
rect 95238 596264 95294 596320
rect 110510 489368 110566 489424
rect 92938 488452 92940 488472
rect 92940 488452 92992 488472
rect 92992 488452 92994 488472
rect 92938 488416 92994 488452
rect 94226 488436 94282 488472
rect 94226 488416 94228 488436
rect 94228 488416 94280 488436
rect 94280 488416 94282 488436
rect 97814 488416 97870 488472
rect 99194 488416 99250 488472
rect 100022 488416 100078 488472
rect 101126 488416 101182 488472
rect 102414 488416 102470 488472
rect 104806 488416 104862 488472
rect 105358 488416 105414 488472
rect 105726 488416 105782 488472
rect 115662 488416 115718 488472
rect 120630 488416 120686 488472
rect 125598 488416 125654 488472
rect 130658 488416 130714 488472
rect 135534 488416 135590 488472
rect 140686 488416 140742 488472
rect 95330 488316 95332 488336
rect 95332 488316 95384 488336
rect 95384 488316 95386 488336
rect 95330 488280 95386 488316
rect 103426 487464 103482 487520
rect 186870 637064 186926 637120
rect 186778 635976 186834 636032
rect 186594 608368 186650 608424
rect 187330 634344 187386 634400
rect 187238 631624 187294 631680
rect 187146 628632 187202 628688
rect 187054 610272 187110 610328
rect 186870 527040 186926 527096
rect 186686 525952 186742 526008
rect 187422 633256 187478 633312
rect 187330 524320 187386 524376
rect 187514 630264 187570 630320
rect 187422 523232 187478 523288
rect 187238 521600 187294 521656
rect 187606 608640 187662 608696
rect 187054 500248 187110 500304
rect 186594 498208 186650 498264
rect 187606 498616 187662 498672
rect 187054 498208 187110 498264
rect 188342 524320 188398 524376
rect 187790 523232 187846 523288
rect 187974 521600 188030 521656
rect 188158 520240 188214 520296
rect 188066 518608 188122 518664
rect 188894 488280 188950 488336
rect 3054 371320 3110 371376
rect 3146 345344 3202 345400
rect 2778 319232 2834 319288
rect 3330 306176 3386 306232
rect 3238 293120 3294 293176
rect 3238 267144 3294 267200
rect 3146 254088 3202 254144
rect 3330 241032 3386 241088
rect 3146 214920 3202 214976
rect 3330 201864 3386 201920
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3146 110608 3202 110664
rect 3238 97552 3294 97608
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 3330 58520 3386 58576
rect 3514 423580 3516 423600
rect 3516 423580 3568 423600
rect 3568 423580 3570 423600
rect 3514 423544 3570 423580
rect 3514 410488 3570 410544
rect 3514 397432 3570 397488
rect 3514 358400 3570 358456
rect 3422 45464 3478 45520
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 570 4800 626 4856
rect 3698 188808 3754 188864
rect 3606 136720 3662 136776
rect 189078 525952 189134 526008
rect 189906 487736 189962 487792
rect 209962 597488 210018 597544
rect 212354 597488 212410 597544
rect 213826 597488 213882 597544
rect 214838 597488 214894 597544
rect 215298 597488 215354 597544
rect 219438 597488 219494 597544
rect 225510 597524 225512 597544
rect 225512 597524 225564 597544
rect 225564 597524 225566 597544
rect 225510 597488 225566 597524
rect 230662 597488 230718 597544
rect 234618 597508 234674 597544
rect 234618 597488 234620 597508
rect 234620 597488 234672 597508
rect 234672 597488 234674 597508
rect 209042 597352 209098 597408
rect 207662 597216 207718 597272
rect 204350 596536 204406 596592
rect 202878 596400 202934 596456
rect 204258 596264 204314 596320
rect 212446 596944 212502 597000
rect 240506 597488 240562 597544
rect 245474 597488 245530 597544
rect 250534 597488 250590 597544
rect 215298 488416 215354 488472
rect 220726 488416 220782 488472
rect 226246 488416 226302 488472
rect 230478 488416 230534 488472
rect 202878 488044 202880 488064
rect 202880 488044 202932 488064
rect 202932 488044 202934 488064
rect 202878 488008 202934 488044
rect 204258 488028 204314 488064
rect 204258 488008 204260 488028
rect 204260 488008 204312 488028
rect 204312 488008 204314 488028
rect 211802 488008 211858 488064
rect 211158 487872 211214 487928
rect 204902 487328 204958 487384
rect 203522 487192 203578 487248
rect 210054 487484 210110 487520
rect 210054 487464 210056 487484
rect 210056 487464 210108 487484
rect 210108 487464 210110 487484
rect 205086 487192 205142 487248
rect 207662 487192 207718 487248
rect 209042 487192 209098 487248
rect 209594 446664 209650 446720
rect 11058 395256 11114 395312
rect 3514 6432 3570 6488
rect 11150 353912 11206 353968
rect 42062 397976 42118 398032
rect 27618 395392 27674 395448
rect 13542 12960 13598 13016
rect 17038 11600 17094 11656
rect 30378 355272 30434 355328
rect 48318 396616 48374 396672
rect 46938 393896 46994 393952
rect 67638 395528 67694 395584
rect 49698 351056 49754 351112
rect 51354 8880 51410 8936
rect 66718 13096 66774 13152
rect 65062 10240 65118 10296
rect 82818 394032 82874 394088
rect 81438 177248 81494 177304
rect 85578 177384 85634 177440
rect 121458 395800 121514 395856
rect 118698 395664 118754 395720
rect 100758 10376 100814 10432
rect 102230 14456 102286 14512
rect 118790 351192 118846 351248
rect 127622 354048 127678 354104
rect 122838 352552 122894 352608
rect 138018 396752 138074 396808
rect 135258 352688 135314 352744
rect 137650 7520 137706 7576
rect 140042 13232 140098 13288
rect 141238 7656 141294 7712
rect 154578 394168 154634 394224
rect 153198 351328 153254 351384
rect 156602 354184 156658 354240
rect 172518 352824 172574 352880
rect 170770 7792 170826 7848
rect 174266 9016 174322 9072
rect 175462 3304 175518 3360
rect 187698 352960 187754 353016
rect 191838 396888 191894 396944
rect 194414 6160 194470 6216
rect 204350 446256 204406 446312
rect 201958 445984 202014 446040
rect 202142 442312 202198 442368
rect 202510 442448 202566 442504
rect 203430 443672 203486 443728
rect 202694 442584 202750 442640
rect 204626 446120 204682 446176
rect 209042 446528 209098 446584
rect 206834 446392 206890 446448
rect 205454 444760 205510 444816
rect 205730 444624 205786 444680
rect 206282 444488 206338 444544
rect 207110 444896 207166 444952
rect 213182 487464 213238 487520
rect 214562 487192 214618 487248
rect 215942 487192 215998 487248
rect 213090 444080 213146 444136
rect 207570 443808 207626 443864
rect 205086 443536 205142 443592
rect 205362 443400 205418 443456
rect 206190 443400 206246 443456
rect 210606 443400 210662 443456
rect 211066 443808 211122 443864
rect 217414 443944 217470 444000
rect 219346 443808 219402 443864
rect 217414 443672 217470 443728
rect 219898 487736 219954 487792
rect 219714 476720 219770 476776
rect 220450 443944 220506 444000
rect 228546 454008 228602 454064
rect 229006 446392 229062 446448
rect 229098 446256 229154 446312
rect 229742 446120 229798 446176
rect 235630 487872 235686 487928
rect 235538 446800 235594 446856
rect 233606 446256 233662 446312
rect 234710 445984 234766 446040
rect 232318 443808 232374 443864
rect 233238 443808 233294 443864
rect 235262 445032 235318 445088
rect 237746 446120 237802 446176
rect 241426 487872 241482 487928
rect 250442 487464 250498 487520
rect 245566 487348 245622 487384
rect 245566 487328 245568 487348
rect 245568 487328 245620 487348
rect 245620 487328 245622 487348
rect 245474 445576 245530 445632
rect 247498 444080 247554 444136
rect 250442 445712 250498 445768
rect 251546 444352 251602 444408
rect 251730 445984 251786 446040
rect 251822 445848 251878 445904
rect 252926 449112 252982 449168
rect 254030 449248 254086 449304
rect 234894 443808 234950 443864
rect 258446 445576 258502 445632
rect 260838 446120 260894 446176
rect 283838 699760 283894 699816
rect 264426 446256 264482 446312
rect 264242 444760 264298 444816
rect 256606 443536 256662 443592
rect 258906 443400 258962 443456
rect 259366 443400 259422 443456
rect 262126 443400 262182 443456
rect 260010 400152 260066 400208
rect 208214 398792 208270 398848
rect 207754 398656 207810 398712
rect 206282 398520 206338 398576
rect 204994 397568 205050 397624
rect 205638 397024 205694 397080
rect 206466 397432 206522 397488
rect 210238 398112 210294 398168
rect 208398 394304 208454 394360
rect 210330 397704 210386 397760
rect 210238 397568 210294 397624
rect 210698 397840 210754 397896
rect 211250 397568 211306 397624
rect 211526 398384 211582 398440
rect 211434 397840 211490 397896
rect 211618 397704 211674 397760
rect 211342 397432 211398 397488
rect 211158 395256 211214 395312
rect 212170 398792 212226 398848
rect 212262 397704 212318 397760
rect 212630 398656 212686 398712
rect 212630 397840 212686 397896
rect 212538 397432 212594 397488
rect 212814 398520 212870 398576
rect 212722 397432 212778 397488
rect 213366 397976 213422 398032
rect 213918 398112 213974 398168
rect 214010 397840 214066 397896
rect 214286 397568 214342 397624
rect 214194 397432 214250 397488
rect 214010 396616 214066 396672
rect 214746 397704 214802 397760
rect 214746 397568 214802 397624
rect 215298 397976 215354 398032
rect 215574 397704 215630 397760
rect 215482 397568 215538 397624
rect 215390 397432 215446 397488
rect 215758 397432 215814 397488
rect 216770 398928 216826 398984
rect 216678 397704 216734 397760
rect 216862 397568 216918 397624
rect 216954 397432 217010 397488
rect 217138 397840 217194 397896
rect 218058 397704 218114 397760
rect 218242 397568 218298 397624
rect 218150 397432 218206 397488
rect 218886 397840 218942 397896
rect 219346 398384 219402 398440
rect 219346 398248 219402 398304
rect 219806 398248 219862 398304
rect 219622 397704 219678 397760
rect 219530 397568 219586 397624
rect 219346 395800 219402 395856
rect 219898 397432 219954 397488
rect 220818 397704 220874 397760
rect 221002 397432 221058 397488
rect 221278 397568 221334 397624
rect 221094 396752 221150 396808
rect 222382 397568 222438 397624
rect 222290 397432 222346 397488
rect 223762 397840 223818 397896
rect 223578 397568 223634 397624
rect 223946 397704 224002 397760
rect 223854 397432 223910 397488
rect 224958 397568 225014 397624
rect 225234 396888 225290 396944
rect 225418 397432 225474 397488
rect 226338 397024 226394 397080
rect 226522 397432 226578 397488
rect 228822 397704 228878 397760
rect 229006 397568 229062 397624
rect 228730 397432 228786 397488
rect 228914 397432 228970 397488
rect 230202 397840 230258 397896
rect 230294 397704 230350 397760
rect 230386 397568 230442 397624
rect 230110 397432 230166 397488
rect 231122 353368 231178 353424
rect 231490 397432 231546 397488
rect 231766 397568 231822 397624
rect 231582 395528 231638 395584
rect 232134 394032 232190 394088
rect 232318 393760 232374 393816
rect 232962 397704 233018 397760
rect 233146 397568 233202 397624
rect 233054 397432 233110 397488
rect 232870 396480 232926 396536
rect 233606 397976 233662 398032
rect 233514 389544 233570 389600
rect 233422 389136 233478 389192
rect 234158 397568 234214 397624
rect 234066 397432 234122 397488
rect 234434 397704 234490 397760
rect 234526 397432 234582 397488
rect 234894 393760 234950 393816
rect 235262 393760 235318 393816
rect 235722 397568 235778 397624
rect 235814 397432 235870 397488
rect 235630 397160 235686 397216
rect 235906 397024 235962 397080
rect 237194 397704 237250 397760
rect 237286 397568 237342 397624
rect 237102 397432 237158 397488
rect 236642 353504 236698 353560
rect 238482 397704 238538 397760
rect 238390 397568 238446 397624
rect 238574 397432 238630 397488
rect 238666 396888 238722 396944
rect 237930 353912 237986 353968
rect 239678 397704 239734 397760
rect 239770 397568 239826 397624
rect 240046 397840 240102 397896
rect 239954 397432 240010 397488
rect 241426 397568 241482 397624
rect 241334 397432 241390 397488
rect 242438 397704 242494 397760
rect 242622 398656 242678 398712
rect 242530 397568 242586 397624
rect 239310 3440 239366 3496
rect 240506 3304 240562 3360
rect 242806 398928 242862 398984
rect 242714 397432 242770 397488
rect 242622 396752 242678 396808
rect 243910 397840 243966 397896
rect 244002 397704 244058 397760
rect 244186 397568 244242 397624
rect 244094 397432 244150 397488
rect 245382 399064 245438 399120
rect 245566 397568 245622 397624
rect 245474 397432 245530 397488
rect 246486 397432 246542 397488
rect 246670 397568 246726 397624
rect 246946 397704 247002 397760
rect 246854 397432 246910 397488
rect 247314 398384 247370 398440
rect 248142 397704 248198 397760
rect 248326 397568 248382 397624
rect 248050 397432 248106 397488
rect 248234 397432 248290 397488
rect 248510 398112 248566 398168
rect 248786 398520 248842 398576
rect 249522 397568 249578 397624
rect 249706 397704 249762 397760
rect 249614 397432 249670 397488
rect 249890 397976 249946 398032
rect 250902 397840 250958 397896
rect 250994 397704 251050 397760
rect 251086 397568 251142 397624
rect 250810 397432 250866 397488
rect 251270 398248 251326 398304
rect 252190 397704 252246 397760
rect 252282 397568 252338 397624
rect 252466 397840 252522 397896
rect 252374 397432 252430 397488
rect 253110 399336 253166 399392
rect 253202 398656 253258 398712
rect 253110 398248 253166 398304
rect 253662 399472 253718 399528
rect 253662 398384 253718 398440
rect 253662 397840 253718 397896
rect 253754 397704 253810 397760
rect 253846 397568 253902 397624
rect 253570 397432 253626 397488
rect 255226 399200 255282 399256
rect 255134 397568 255190 397624
rect 255042 397432 255098 397488
rect 254674 5344 254730 5400
rect 257250 399064 257306 399120
rect 257250 398656 257306 398712
rect 255594 398248 255650 398304
rect 255594 395664 255650 395720
rect 256238 398520 256294 398576
rect 256790 398248 256846 398304
rect 258814 398520 258870 398576
rect 263506 398656 263562 398712
rect 261482 397704 261538 397760
rect 258262 5208 258318 5264
rect 263414 398384 263470 398440
rect 265806 445848 265862 445904
rect 265714 444624 265770 444680
rect 265622 443536 265678 443592
rect 267002 444488 267058 444544
rect 281814 596808 281870 596864
rect 284666 597216 284722 597272
rect 284390 596944 284446 597000
rect 284758 597080 284814 597136
rect 282366 488008 282422 488064
rect 284666 449248 284722 449304
rect 285586 489776 285642 489832
rect 285034 488552 285090 488608
rect 285586 488552 285642 488608
rect 298006 636928 298062 636984
rect 297914 635840 297970 635896
rect 297822 634208 297878 634264
rect 297638 633120 297694 633176
rect 297454 631488 297510 631544
rect 296994 610136 297050 610192
rect 296902 608232 296958 608288
rect 297086 608640 297142 608696
rect 296994 500792 297050 500848
rect 297546 628496 297602 628552
rect 297454 521600 297510 521656
rect 297730 630128 297786 630184
rect 297730 527040 297786 527096
rect 298006 525972 298062 526008
rect 298006 525952 298008 525972
rect 298008 525952 298060 525972
rect 298060 525952 298062 525972
rect 298006 524320 298062 524376
rect 297914 523232 297970 523288
rect 297822 520240 297878 520296
rect 297546 518608 297602 518664
rect 297914 500792 297970 500848
rect 297914 500248 297970 500304
rect 297454 498616 297510 498672
rect 296902 498208 296958 498264
rect 284758 449112 284814 449168
rect 297822 498208 297878 498264
rect 319994 597488 320050 597544
rect 322294 597488 322350 597544
rect 323398 597488 323454 597544
rect 324778 597488 324834 597544
rect 326158 597508 326214 597544
rect 326158 597488 326160 597508
rect 326160 597488 326212 597508
rect 326212 597488 326214 597508
rect 314658 597352 314714 597408
rect 330390 597488 330446 597544
rect 335358 597524 335360 597544
rect 335360 597524 335412 597544
rect 335412 597524 335414 597544
rect 335358 597488 335414 597524
rect 340510 597488 340566 597544
rect 345662 597488 345718 597544
rect 350446 597488 350502 597544
rect 354678 597488 354734 597544
rect 360566 597488 360622 597544
rect 311898 596284 311954 596320
rect 311898 596264 311900 596284
rect 311900 596264 311952 596284
rect 311952 596264 311954 596284
rect 313278 596264 313334 596320
rect 325330 489096 325386 489152
rect 330482 488416 330538 488472
rect 335450 488416 335506 488472
rect 340602 488452 340604 488472
rect 340604 488452 340656 488472
rect 340656 488452 340658 488472
rect 340602 488416 340658 488452
rect 345754 488416 345810 488472
rect 350354 488416 350410 488472
rect 355782 488416 355838 488472
rect 360474 488416 360530 488472
rect 313922 488280 313978 488336
rect 312542 487192 312598 487248
rect 315302 488144 315358 488200
rect 318890 487872 318946 487928
rect 318062 487192 318118 487248
rect 323582 487328 323638 487384
rect 319442 487192 319498 487248
rect 320086 487192 320142 487248
rect 320822 487192 320878 487248
rect 322202 487192 322258 487248
rect 324870 487212 324926 487248
rect 324870 487192 324872 487212
rect 324872 487192 324924 487212
rect 324924 487192 324926 487212
rect 326342 487192 326398 487248
rect 407762 636384 407818 636440
rect 407578 630944 407634 631000
rect 407394 627952 407450 628008
rect 407946 635296 408002 635352
rect 407854 607688 407910 607744
rect 407486 527040 407542 527096
rect 407670 526496 407726 526552
rect 407670 523232 407726 523288
rect 407578 520920 407634 520976
rect 407486 517928 407542 517984
rect 408222 633664 408278 633720
rect 408038 632576 408094 632632
rect 407854 498344 407910 498400
rect 408130 629584 408186 629640
rect 408038 523232 408094 523288
rect 408406 610000 408462 610056
rect 408314 608640 408370 608696
rect 408130 520240 408186 520296
rect 408038 498208 408094 498264
rect 407946 488280 408002 488336
rect 407762 488144 407818 488200
rect 407486 488008 407542 488064
rect 408406 500248 408462 500304
rect 408314 498616 408370 498672
rect 408314 498208 408370 498264
rect 429198 597488 429254 597544
rect 434718 597508 434774 597544
rect 434718 597488 434720 597508
rect 434720 597488 434772 597508
rect 434772 597488 434774 597508
rect 444378 597524 444380 597544
rect 444380 597524 444432 597544
rect 444432 597524 444434 597544
rect 444378 597488 444434 597524
rect 459558 597488 459614 597544
rect 440238 597372 440294 597408
rect 440238 597352 440240 597372
rect 440240 597352 440292 597372
rect 440292 597352 440294 597372
rect 455418 597352 455474 597408
rect 465078 597352 465134 597408
rect 433338 597216 433394 597272
rect 449898 597236 449954 597272
rect 449898 597216 449900 597236
rect 449900 597216 449952 597236
rect 449952 597216 449954 597236
rect 434718 597100 434774 597136
rect 434718 597080 434720 597100
rect 434720 597080 434772 597100
rect 434772 597080 434774 597100
rect 431958 596828 432014 596864
rect 431958 596808 431960 596828
rect 431960 596808 432012 596828
rect 432012 596808 432014 596828
rect 470598 596964 470654 597000
rect 470598 596944 470600 596964
rect 470600 596944 470652 596964
rect 470652 596944 470654 596964
rect 422574 596400 422630 596456
rect 423678 596284 423734 596320
rect 423678 596264 423680 596284
rect 423680 596264 423732 596284
rect 423732 596264 423734 596284
rect 425058 596264 425114 596320
rect 422574 488436 422630 488472
rect 422574 488416 422576 488436
rect 422576 488416 422628 488436
rect 422628 488416 422630 488436
rect 423678 488452 423680 488472
rect 423680 488452 423732 488472
rect 423732 488452 423734 488472
rect 423678 488416 423734 488452
rect 434718 488416 434774 488472
rect 440238 488416 440294 488472
rect 444378 488416 444434 488472
rect 449898 488416 449954 488472
rect 430578 488280 430634 488336
rect 465078 488280 465134 488336
rect 427818 488164 427874 488200
rect 427818 488144 427820 488164
rect 427820 488144 427872 488164
rect 427872 488144 427874 488164
rect 429198 488144 429254 488200
rect 426438 487756 426494 487792
rect 426438 487736 426440 487756
rect 426440 487736 426492 487756
rect 426492 487736 426494 487756
rect 434718 488144 434774 488200
rect 455418 488008 455474 488064
rect 459558 487872 459614 487928
rect 470598 488028 470654 488064
rect 470598 488008 470600 488028
rect 470600 488008 470652 488028
rect 470652 488008 470654 488028
rect 432050 487600 432106 487656
rect 433338 487328 433394 487384
rect 434718 487212 434774 487248
rect 434718 487192 434720 487212
rect 434720 487192 434772 487212
rect 434772 487192 434774 487212
rect 298006 452376 298062 452432
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580262 577632 580318 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 297362 448296 297418 448352
rect 298926 446528 298982 446584
rect 296074 445984 296130 446040
rect 272522 444896 272578 444952
rect 295982 443128 296038 443184
rect 273258 395528 273314 395584
rect 272430 9016 272486 9072
rect 276110 17448 276166 17504
rect 289818 396480 289874 396536
rect 291198 87624 291254 87680
rect 292578 18536 292634 18592
rect 296166 443264 296222 443320
rect 296626 442176 296682 442232
rect 296994 404096 297050 404152
rect 298006 443536 298062 443592
rect 298006 439456 298062 439512
rect 298006 434696 298062 434752
rect 298006 430616 298062 430672
rect 298006 425856 298062 425912
rect 297914 421776 297970 421832
rect 297638 417016 297694 417072
rect 297546 412936 297602 412992
rect 298006 408176 298062 408232
rect 298742 443672 298798 443728
rect 383934 454008 383990 454064
rect 384026 452240 384082 452296
rect 384026 448160 384082 448216
rect 383934 438640 383990 438696
rect 383934 421640 383990 421696
rect 385498 442856 385554 442912
rect 385406 434016 385462 434072
rect 580170 431568 580226 431624
rect 385314 429936 385370 429992
rect 385222 425176 385278 425232
rect 580262 418240 580318 418296
rect 385130 416336 385186 416392
rect 385038 412256 385094 412312
rect 385038 407496 385094 407552
rect 579986 404912 580042 404968
rect 312266 399064 312322 399120
rect 324502 399064 324558 399120
rect 316130 398248 316186 398304
rect 310518 397296 310574 397352
rect 292578 7792 292634 7848
rect 304998 354320 305054 354376
rect 299662 3712 299718 3768
rect 306746 7656 306802 7712
rect 324318 397160 324374 397216
rect 310242 7520 310298 7576
rect 328458 397024 328514 397080
rect 325698 393896 325754 393952
rect 327998 8880 328054 8936
rect 332874 398384 332930 398440
rect 379242 398792 379298 398848
rect 362498 398656 362554 398712
rect 357990 398520 358046 398576
rect 580262 399472 580318 399528
rect 364338 396888 364394 396944
rect 345018 355544 345074 355600
rect 343638 25472 343694 25528
rect 346398 352960 346454 353016
rect 360198 355408 360254 355464
rect 363510 10512 363566 10568
rect 362314 5072 362370 5128
rect 378138 20168 378194 20224
rect 377678 10376 377734 10432
rect 381174 10240 381230 10296
rect 382370 20032 382426 20088
rect 398838 351192 398894 351248
rect 416778 396752 416834 396808
rect 414018 352824 414074 352880
rect 398930 11872 398986 11928
rect 412638 11736 412694 11792
rect 431958 354184 432014 354240
rect 415490 11600 415546 11656
rect 432050 87488 432106 87544
rect 434718 21256 434774 21312
rect 433982 13096 434038 13152
rect 452658 354048 452714 354104
rect 451646 12960 451702 13016
rect 489918 398112 489974 398168
rect 465078 26832 465134 26888
rect 466458 22752 466514 22808
rect 470598 19896 470654 19952
rect 469862 14728 469918 14784
rect 485778 352688 485834 352744
rect 484766 14592 484822 14648
rect 488814 14456 488870 14512
rect 487618 3576 487674 3632
rect 507858 397976 507914 398032
rect 506478 355272 506534 355328
rect 503718 22616 503774 22672
rect 505374 4936 505430 4992
rect 521658 395392 521714 395448
rect 520278 15952 520334 16008
rect 523774 15816 523830 15872
rect 523038 3440 523094 3496
rect 540978 352552 541034 352608
rect 538218 351056 538274 351112
rect 539598 24248 539654 24304
rect 540794 4800 540850 4856
rect 556158 395256 556214 395312
rect 557538 353912 557594 353968
rect 556250 17312 556306 17368
rect 558918 17176 558974 17232
rect 576858 396616 576914 396672
rect 574098 24112 574154 24168
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580170 165824 580226 165880
rect 580262 152632 580318 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 576306 6160 576362 6216
rect 580262 6568 580318 6624
rect 579802 3304 579858 3360
<< metal3 >>
rect 282126 699756 282132 699820
rect 282196 699818 282202 699820
rect 283833 699818 283899 699821
rect 282196 699816 283899 699818
rect 282196 699760 283838 699816
rect 283894 699760 283899 699816
rect 282196 699758 283899 699760
rect 282196 699756 282202 699758
rect 283833 699755 283899 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 186865 637122 186931 637125
rect 186865 637120 189458 637122
rect 186865 637064 186870 637120
rect 186926 637064 189458 637120
rect 186865 637062 189458 637064
rect 186865 637059 186931 637062
rect 189398 637060 189458 637062
rect 78581 636442 78647 636445
rect 80002 636442 80062 637030
rect 189398 637000 190072 637060
rect 299430 637000 300012 637060
rect 298001 636986 298067 636989
rect 299430 636986 299490 637000
rect 298001 636984 299490 636986
rect 298001 636928 298006 636984
rect 298062 636928 299490 636984
rect 298001 636926 299490 636928
rect 298001 636923 298067 636926
rect 78581 636440 80062 636442
rect 78581 636384 78586 636440
rect 78642 636384 80062 636440
rect 78581 636382 80062 636384
rect 407757 636442 407823 636445
rect 410002 636442 410062 637030
rect 407757 636440 410062 636442
rect 407757 636384 407762 636440
rect 407818 636384 410062 636440
rect 407757 636382 410062 636384
rect 78581 636379 78647 636382
rect 407757 636379 407823 636382
rect 186773 636034 186839 636037
rect 186773 636032 189458 636034
rect 186773 635976 186778 636032
rect 186834 635976 189458 636032
rect 186773 635974 189458 635976
rect 186773 635971 186839 635974
rect 189398 635972 189458 635974
rect 78305 635354 78371 635357
rect 80002 635354 80062 635942
rect 189398 635912 190072 635972
rect 299430 635912 300012 635972
rect 297909 635898 297975 635901
rect 299430 635898 299490 635912
rect 297909 635896 299490 635898
rect 297909 635840 297914 635896
rect 297970 635840 299490 635896
rect 297909 635838 299490 635840
rect 297909 635835 297975 635838
rect 78305 635352 80062 635354
rect 78305 635296 78310 635352
rect 78366 635296 80062 635352
rect 78305 635294 80062 635296
rect 407941 635354 408007 635357
rect 410002 635354 410062 635942
rect 407941 635352 410062 635354
rect 407941 635296 407946 635352
rect 408002 635296 410062 635352
rect 407941 635294 410062 635296
rect 78305 635291 78371 635294
rect 407941 635291 408007 635294
rect 187325 634402 187391 634405
rect 187325 634400 189458 634402
rect 187325 634344 187330 634400
rect 187386 634344 189458 634400
rect 187325 634342 189458 634344
rect 187325 634339 187391 634342
rect 189398 634340 189458 634342
rect 78213 633722 78279 633725
rect 80002 633722 80062 634310
rect 189398 634280 190072 634340
rect 299430 634280 300012 634340
rect 297817 634266 297883 634269
rect 299430 634266 299490 634280
rect 297817 634264 299490 634266
rect 297817 634208 297822 634264
rect 297878 634208 299490 634264
rect 297817 634206 299490 634208
rect 297817 634203 297883 634206
rect 78213 633720 80062 633722
rect 78213 633664 78218 633720
rect 78274 633664 80062 633720
rect 78213 633662 80062 633664
rect 408217 633722 408283 633725
rect 410002 633722 410062 634310
rect 408217 633720 410062 633722
rect 408217 633664 408222 633720
rect 408278 633664 410062 633720
rect 408217 633662 410062 633664
rect 78213 633659 78279 633662
rect 408217 633659 408283 633662
rect 187417 633314 187483 633317
rect 187417 633312 189458 633314
rect 187417 633256 187422 633312
rect 187478 633256 189458 633312
rect 187417 633254 189458 633256
rect 187417 633251 187483 633254
rect 189398 633252 189458 633254
rect 77937 632634 78003 632637
rect 80002 632634 80062 633222
rect 189398 633192 190072 633252
rect 299430 633192 300012 633252
rect 297633 633178 297699 633181
rect 299430 633178 299490 633192
rect 297633 633176 299490 633178
rect 297633 633120 297638 633176
rect 297694 633120 299490 633176
rect 297633 633118 299490 633120
rect 297633 633115 297699 633118
rect 77937 632632 80062 632634
rect 77937 632576 77942 632632
rect 77998 632576 80062 632632
rect 77937 632574 80062 632576
rect 408033 632634 408099 632637
rect 410002 632634 410062 633222
rect 408033 632632 410062 632634
rect 408033 632576 408038 632632
rect 408094 632576 410062 632632
rect 408033 632574 410062 632576
rect 77937 632571 78003 632574
rect 408033 632571 408099 632574
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 187233 631682 187299 631685
rect 187233 631680 189458 631682
rect 187233 631624 187238 631680
rect 187294 631624 189458 631680
rect 187233 631622 189458 631624
rect 187233 631619 187299 631622
rect 189398 631620 189458 631622
rect 78121 631002 78187 631005
rect 80002 631002 80062 631590
rect 189398 631560 190072 631620
rect 299430 631560 300012 631620
rect 297449 631546 297515 631549
rect 299430 631546 299490 631560
rect 297449 631544 299490 631546
rect 297449 631488 297454 631544
rect 297510 631488 299490 631544
rect 297449 631486 299490 631488
rect 297449 631483 297515 631486
rect 78121 631000 80062 631002
rect 78121 630944 78126 631000
rect 78182 630944 80062 631000
rect 78121 630942 80062 630944
rect 407573 631002 407639 631005
rect 410002 631002 410062 631590
rect 407573 631000 410062 631002
rect 407573 630944 407578 631000
rect 407634 630944 410062 631000
rect 407573 630942 410062 630944
rect 78121 630939 78187 630942
rect 407573 630939 407639 630942
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 187509 630322 187575 630325
rect 187509 630320 189458 630322
rect 187509 630264 187514 630320
rect 187570 630264 189458 630320
rect 187509 630262 189458 630264
rect 187509 630259 187575 630262
rect 189398 630260 189458 630262
rect 77753 629642 77819 629645
rect 80002 629642 80062 630230
rect 189398 630200 190072 630260
rect 299430 630200 300012 630260
rect 297725 630186 297791 630189
rect 299430 630186 299490 630200
rect 297725 630184 299490 630186
rect 297725 630128 297730 630184
rect 297786 630128 299490 630184
rect 297725 630126 299490 630128
rect 297725 630123 297791 630126
rect 77753 629640 80062 629642
rect 77753 629584 77758 629640
rect 77814 629584 80062 629640
rect 77753 629582 80062 629584
rect 408125 629642 408191 629645
rect 410002 629642 410062 630230
rect 408125 629640 410062 629642
rect 408125 629584 408130 629640
rect 408186 629584 410062 629640
rect 408125 629582 410062 629584
rect 77753 629579 77819 629582
rect 408125 629579 408191 629582
rect 187141 628690 187207 628693
rect 187141 628688 189458 628690
rect 187141 628632 187146 628688
rect 187202 628632 189458 628688
rect 187141 628630 189458 628632
rect 187141 628627 187207 628630
rect 189398 628628 189458 628630
rect 78029 628010 78095 628013
rect 80002 628010 80062 628598
rect 189398 628568 190072 628628
rect 299430 628568 300012 628628
rect 297541 628554 297607 628557
rect 299430 628554 299490 628568
rect 297541 628552 299490 628554
rect 297541 628496 297546 628552
rect 297602 628496 299490 628552
rect 297541 628494 299490 628496
rect 297541 628491 297607 628494
rect 78029 628008 80062 628010
rect 78029 627952 78034 628008
rect 78090 627952 80062 628008
rect 78029 627950 80062 627952
rect 407389 628010 407455 628013
rect 410002 628010 410062 628598
rect 407389 628008 410062 628010
rect 407389 627952 407394 628008
rect 407450 627952 410062 628008
rect 407389 627950 410062 627952
rect 78029 627947 78095 627950
rect 407389 627947 407455 627950
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 187049 610330 187115 610333
rect 187049 610328 189458 610330
rect 187049 610272 187054 610328
rect 187110 610272 189458 610328
rect 187049 610270 189458 610272
rect 187049 610267 187115 610270
rect 189398 610268 189458 610270
rect 78397 610058 78463 610061
rect 80002 610058 80062 610238
rect 189398 610208 190072 610268
rect 299430 610208 300012 610268
rect 296989 610194 297055 610197
rect 299430 610194 299490 610208
rect 296989 610192 299490 610194
rect 296989 610136 296994 610192
rect 297050 610136 299490 610192
rect 296989 610134 299490 610136
rect 296989 610131 297055 610134
rect 78397 610056 80062 610058
rect 78397 610000 78402 610056
rect 78458 610000 80062 610056
rect 78397 609998 80062 610000
rect 408401 610058 408467 610061
rect 410002 610058 410062 610238
rect 408401 610056 410062 610058
rect 408401 610000 408406 610056
rect 408462 610000 410062 610056
rect 408401 609998 410062 610000
rect 78397 609995 78463 609998
rect 408401 609995 408467 609998
rect 77845 608698 77911 608701
rect 187601 608698 187667 608701
rect 297081 608698 297147 608701
rect 408309 608698 408375 608701
rect 77845 608696 80062 608698
rect 77845 608640 77850 608696
rect 77906 608640 80062 608696
rect 77845 608638 80062 608640
rect 77845 608635 77911 608638
rect 80002 608606 80062 608638
rect 187601 608696 189458 608698
rect 187601 608640 187606 608696
rect 187662 608640 189458 608696
rect 187601 608638 189458 608640
rect 187601 608635 187667 608638
rect 189398 608636 189458 608638
rect 297081 608696 299490 608698
rect 297081 608640 297086 608696
rect 297142 608640 299490 608696
rect 297081 608638 299490 608640
rect 189398 608576 190072 608636
rect 297081 608635 297147 608638
rect 299430 608636 299490 608638
rect 408309 608696 410062 608698
rect 408309 608640 408314 608696
rect 408370 608640 410062 608696
rect 408309 608638 410062 608640
rect 299430 608576 300012 608636
rect 408309 608635 408375 608638
rect 410002 608606 410062 608638
rect 186589 608426 186655 608429
rect 186589 608424 189458 608426
rect 186589 608368 186594 608424
rect 186650 608368 189458 608424
rect 186589 608366 189458 608368
rect 186589 608363 186655 608366
rect 189398 608364 189458 608366
rect 78581 607746 78647 607749
rect 80002 607746 80062 608334
rect 189398 608304 190072 608364
rect 299430 608304 300012 608364
rect 296897 608290 296963 608293
rect 299430 608290 299490 608304
rect 296897 608288 299490 608290
rect 296897 608232 296902 608288
rect 296958 608232 299490 608288
rect 296897 608230 299490 608232
rect 296897 608227 296963 608230
rect 78581 607744 80062 607746
rect 78581 607688 78586 607744
rect 78642 607688 80062 607744
rect 78581 607686 80062 607688
rect 407849 607746 407915 607749
rect 410002 607746 410062 608334
rect 407849 607744 410062 607746
rect 407849 607688 407854 607744
rect 407910 607688 410062 607744
rect 407849 607686 410062 607688
rect 78581 607683 78647 607686
rect 407849 607683 407915 607686
rect -960 606114 480 606204
rect 3141 606114 3207 606117
rect -960 606112 3207 606114
rect -960 606056 3146 606112
rect 3202 606056 3207 606112
rect -960 606054 3207 606056
rect -960 605964 480 606054
rect 3141 606051 3207 606054
rect 583520 604060 584960 604300
rect 102358 597484 102364 597548
rect 102428 597546 102434 597548
rect 103145 597546 103211 597549
rect 102428 597544 103211 597546
rect 102428 597488 103150 597544
rect 103206 597488 103211 597544
rect 102428 597486 103211 597488
rect 102428 597484 102434 597486
rect 103145 597483 103211 597486
rect 105302 597484 105308 597548
rect 105372 597546 105378 597548
rect 106222 597546 106228 597548
rect 105372 597486 106228 597546
rect 105372 597484 105378 597486
rect 106222 597484 106228 597486
rect 106292 597484 106298 597548
rect 110454 597484 110460 597548
rect 110524 597546 110530 597548
rect 111701 597546 111767 597549
rect 110524 597544 111767 597546
rect 110524 597488 111706 597544
rect 111762 597488 111767 597544
rect 110524 597486 111767 597488
rect 110524 597484 110530 597486
rect 111701 597483 111767 597486
rect 115606 597484 115612 597548
rect 115676 597546 115682 597548
rect 115841 597546 115907 597549
rect 115676 597544 115907 597546
rect 115676 597488 115846 597544
rect 115902 597488 115907 597544
rect 115676 597486 115907 597488
rect 115676 597484 115682 597486
rect 115841 597483 115907 597486
rect 120574 597484 120580 597548
rect 120644 597546 120650 597548
rect 121361 597546 121427 597549
rect 120644 597544 121427 597546
rect 120644 597488 121366 597544
rect 121422 597488 121427 597544
rect 120644 597486 121427 597488
rect 120644 597484 120650 597486
rect 121361 597483 121427 597486
rect 125542 597484 125548 597548
rect 125612 597546 125618 597548
rect 126881 597546 126947 597549
rect 125612 597544 126947 597546
rect 125612 597488 126886 597544
rect 126942 597488 126947 597544
rect 125612 597486 126947 597488
rect 125612 597484 125618 597486
rect 126881 597483 126947 597486
rect 130510 597484 130516 597548
rect 130580 597546 130586 597548
rect 131021 597546 131087 597549
rect 130580 597544 131087 597546
rect 130580 597488 131026 597544
rect 131082 597488 131087 597544
rect 130580 597486 131087 597488
rect 130580 597484 130586 597486
rect 131021 597483 131087 597486
rect 135478 597484 135484 597548
rect 135548 597546 135554 597548
rect 136541 597546 136607 597549
rect 140681 597548 140747 597549
rect 135548 597544 136607 597546
rect 135548 597488 136546 597544
rect 136602 597488 136607 597544
rect 135548 597486 136607 597488
rect 135548 597484 135554 597486
rect 136541 597483 136607 597486
rect 140630 597484 140636 597548
rect 140700 597546 140747 597548
rect 209957 597548 210023 597549
rect 212349 597548 212415 597549
rect 140700 597544 140792 597546
rect 140742 597488 140792 597544
rect 140700 597486 140792 597488
rect 209957 597544 210004 597548
rect 210068 597546 210074 597548
rect 209957 597488 209962 597544
rect 140700 597484 140747 597486
rect 140681 597483 140747 597484
rect 209957 597484 210004 597488
rect 210068 597486 210114 597546
rect 212349 597544 212396 597548
rect 212460 597546 212466 597548
rect 212349 597488 212354 597544
rect 210068 597484 210074 597486
rect 212349 597484 212396 597488
rect 212460 597486 212506 597546
rect 212460 597484 212466 597486
rect 213494 597484 213500 597548
rect 213564 597546 213570 597548
rect 213821 597546 213887 597549
rect 214833 597548 214899 597549
rect 214782 597546 214788 597548
rect 213564 597544 213887 597546
rect 213564 597488 213826 597544
rect 213882 597488 213887 597544
rect 213564 597486 213887 597488
rect 214742 597486 214788 597546
rect 214852 597544 214899 597548
rect 214894 597488 214899 597544
rect 213564 597484 213570 597486
rect 209957 597483 210023 597484
rect 212349 597483 212415 597484
rect 213821 597483 213887 597486
rect 214782 597484 214788 597486
rect 214852 597484 214899 597488
rect 214833 597483 214899 597484
rect 215293 597546 215359 597549
rect 215702 597546 215708 597548
rect 215293 597544 215708 597546
rect 215293 597488 215298 597544
rect 215354 597488 215708 597544
rect 215293 597486 215708 597488
rect 215293 597483 215359 597486
rect 215702 597484 215708 597486
rect 215772 597484 215778 597548
rect 219198 597484 219204 597548
rect 219268 597546 219274 597548
rect 219433 597546 219499 597549
rect 225505 597548 225571 597549
rect 230657 597548 230723 597549
rect 225454 597546 225460 597548
rect 219268 597544 219499 597546
rect 219268 597488 219438 597544
rect 219494 597488 219499 597544
rect 219268 597486 219499 597488
rect 225414 597486 225460 597546
rect 225524 597544 225571 597548
rect 230606 597546 230612 597548
rect 225566 597488 225571 597544
rect 219268 597484 219274 597486
rect 219433 597483 219499 597486
rect 225454 597484 225460 597486
rect 225524 597484 225571 597488
rect 230566 597486 230612 597546
rect 230676 597544 230723 597548
rect 230718 597488 230723 597544
rect 230606 597484 230612 597486
rect 230676 597484 230723 597488
rect 225505 597483 225571 597484
rect 230657 597483 230723 597484
rect 234613 597546 234679 597549
rect 240501 597548 240567 597549
rect 245469 597548 245535 597549
rect 250529 597548 250595 597549
rect 235574 597546 235580 597548
rect 234613 597544 235580 597546
rect 234613 597488 234618 597544
rect 234674 597488 235580 597544
rect 234613 597486 235580 597488
rect 234613 597483 234679 597486
rect 235574 597484 235580 597486
rect 235644 597484 235650 597548
rect 240501 597544 240548 597548
rect 240612 597546 240618 597548
rect 240501 597488 240506 597544
rect 240501 597484 240548 597488
rect 240612 597486 240658 597546
rect 245469 597544 245516 597548
rect 245580 597546 245586 597548
rect 250478 597546 250484 597548
rect 245469 597488 245474 597544
rect 240612 597484 240618 597486
rect 245469 597484 245516 597488
rect 245580 597486 245626 597546
rect 250438 597486 250484 597546
rect 250548 597544 250595 597548
rect 250590 597488 250595 597544
rect 245580 597484 245586 597486
rect 250478 597484 250484 597486
rect 250548 597484 250595 597488
rect 240501 597483 240567 597484
rect 245469 597483 245535 597484
rect 250529 597483 250595 597484
rect 319989 597548 320055 597549
rect 322289 597548 322355 597549
rect 323393 597548 323459 597549
rect 319989 597544 320036 597548
rect 320100 597546 320106 597548
rect 322238 597546 322244 597548
rect 319989 597488 319994 597544
rect 319989 597484 320036 597488
rect 320100 597486 320146 597546
rect 322198 597486 322244 597546
rect 322308 597544 322355 597548
rect 323342 597546 323348 597548
rect 322350 597488 322355 597544
rect 320100 597484 320106 597486
rect 322238 597484 322244 597486
rect 322308 597484 322355 597488
rect 323302 597486 323348 597546
rect 323412 597544 323459 597548
rect 323454 597488 323459 597544
rect 323342 597484 323348 597486
rect 323412 597484 323459 597488
rect 319989 597483 320055 597484
rect 322289 597483 322355 597484
rect 323393 597483 323459 597484
rect 324773 597548 324839 597549
rect 324773 597544 324820 597548
rect 324884 597546 324890 597548
rect 324773 597488 324778 597544
rect 324773 597484 324820 597488
rect 324884 597486 324930 597546
rect 324884 597484 324890 597486
rect 325734 597484 325740 597548
rect 325804 597546 325810 597548
rect 326153 597546 326219 597549
rect 325804 597544 326219 597546
rect 325804 597488 326158 597544
rect 326214 597488 326219 597544
rect 325804 597486 326219 597488
rect 325804 597484 325810 597486
rect 324773 597483 324839 597484
rect 326153 597483 326219 597486
rect 330385 597546 330451 597549
rect 330518 597546 330524 597548
rect 330385 597544 330524 597546
rect 330385 597488 330390 597544
rect 330446 597488 330524 597544
rect 330385 597486 330524 597488
rect 330385 597483 330451 597486
rect 330518 597484 330524 597486
rect 330588 597484 330594 597548
rect 335118 597484 335124 597548
rect 335188 597546 335194 597548
rect 335353 597546 335419 597549
rect 340505 597548 340571 597549
rect 345657 597548 345723 597549
rect 350441 597548 350507 597549
rect 340454 597546 340460 597548
rect 335188 597544 335419 597546
rect 335188 597488 335358 597544
rect 335414 597488 335419 597544
rect 335188 597486 335419 597488
rect 340414 597486 340460 597546
rect 340524 597544 340571 597548
rect 345606 597546 345612 597548
rect 340566 597488 340571 597544
rect 335188 597484 335194 597486
rect 335353 597483 335419 597486
rect 340454 597484 340460 597486
rect 340524 597484 340571 597488
rect 345566 597486 345612 597546
rect 345676 597544 345723 597548
rect 350390 597546 350396 597548
rect 345718 597488 345723 597544
rect 345606 597484 345612 597486
rect 345676 597484 345723 597488
rect 350350 597486 350396 597546
rect 350460 597544 350507 597548
rect 350502 597488 350507 597544
rect 350390 597484 350396 597486
rect 350460 597484 350507 597488
rect 354438 597484 354444 597548
rect 354508 597546 354514 597548
rect 354673 597546 354739 597549
rect 360561 597548 360627 597549
rect 360510 597546 360516 597548
rect 354508 597544 354739 597546
rect 354508 597488 354678 597544
rect 354734 597488 354739 597544
rect 354508 597486 354739 597488
rect 360470 597486 360516 597546
rect 360580 597544 360627 597548
rect 360622 597488 360627 597544
rect 354508 597484 354514 597486
rect 340505 597483 340571 597484
rect 345657 597483 345723 597484
rect 350441 597483 350507 597484
rect 354673 597483 354739 597486
rect 360510 597484 360516 597486
rect 360580 597484 360627 597488
rect 360561 597483 360627 597484
rect 429193 597546 429259 597549
rect 429878 597546 429884 597548
rect 429193 597544 429884 597546
rect 429193 597488 429198 597544
rect 429254 597488 429884 597544
rect 429193 597486 429884 597488
rect 429193 597483 429259 597486
rect 429878 597484 429884 597486
rect 429948 597484 429954 597548
rect 434713 597546 434779 597549
rect 435582 597546 435588 597548
rect 434713 597544 435588 597546
rect 434713 597488 434718 597544
rect 434774 597488 435588 597544
rect 434713 597486 435588 597488
rect 434713 597483 434779 597486
rect 435582 597484 435588 597486
rect 435652 597484 435658 597548
rect 444373 597546 444439 597549
rect 445518 597546 445524 597548
rect 444373 597544 445524 597546
rect 444373 597488 444378 597544
rect 444434 597488 445524 597544
rect 444373 597486 445524 597488
rect 444373 597483 444439 597486
rect 445518 597484 445524 597486
rect 445588 597484 445594 597548
rect 459553 597546 459619 597549
rect 460422 597546 460428 597548
rect 459553 597544 460428 597546
rect 459553 597488 459558 597544
rect 459614 597488 460428 597544
rect 459553 597486 460428 597488
rect 459553 597483 459619 597486
rect 460422 597484 460428 597486
rect 460492 597484 460498 597548
rect 92473 597410 92539 597413
rect 92974 597410 92980 597412
rect 92473 597408 92980 597410
rect 92473 597352 92478 597408
rect 92534 597352 92980 597408
rect 92473 597350 92980 597352
rect 92473 597347 92539 597350
rect 92974 597348 92980 597350
rect 93044 597348 93050 597412
rect 98862 597348 98868 597412
rect 98932 597410 98938 597412
rect 208894 597410 208900 597412
rect 98932 597350 208900 597410
rect 98932 597348 98938 597350
rect 208894 597348 208900 597350
rect 208964 597410 208970 597412
rect 209037 597410 209103 597413
rect 208964 597408 209103 597410
rect 208964 597352 209042 597408
rect 209098 597352 209103 597408
rect 208964 597350 209103 597352
rect 208964 597348 208970 597350
rect 209037 597347 209103 597350
rect 314653 597410 314719 597413
rect 315246 597410 315252 597412
rect 314653 597408 315252 597410
rect 314653 597352 314658 597408
rect 314714 597352 315252 597408
rect 314653 597350 315252 597352
rect 314653 597347 314719 597350
rect 315246 597348 315252 597350
rect 315316 597348 315322 597412
rect 321134 597348 321140 597412
rect 321204 597410 321210 597412
rect 430982 597410 430988 597412
rect 321204 597350 430988 597410
rect 321204 597348 321210 597350
rect 430982 597348 430988 597350
rect 431052 597348 431058 597412
rect 440233 597410 440299 597413
rect 455413 597412 455479 597413
rect 440366 597410 440372 597412
rect 440233 597408 440372 597410
rect 440233 597352 440238 597408
rect 440294 597352 440372 597408
rect 440233 597350 440372 597352
rect 440233 597347 440299 597350
rect 440366 597348 440372 597350
rect 440436 597348 440442 597412
rect 455413 597410 455460 597412
rect 455368 597408 455460 597410
rect 455368 597352 455418 597408
rect 455368 597350 455460 597352
rect 455413 597348 455460 597350
rect 455524 597348 455530 597412
rect 465073 597410 465139 597413
rect 465390 597410 465396 597412
rect 465073 597408 465396 597410
rect 465073 597352 465078 597408
rect 465134 597352 465396 597408
rect 465073 597350 465396 597352
rect 455413 597347 455479 597348
rect 465073 597347 465139 597350
rect 465390 597348 465396 597350
rect 465460 597348 465466 597412
rect 207657 597276 207723 597277
rect 97758 597212 97764 597276
rect 97828 597274 97834 597276
rect 207606 597274 207612 597276
rect 97828 597214 207612 597274
rect 207676 597274 207723 597276
rect 284661 597274 284727 597277
rect 433333 597276 433399 597277
rect 318926 597274 318932 597276
rect 207676 597272 207804 597274
rect 207718 597216 207804 597272
rect 97828 597212 97834 597214
rect 207606 597212 207612 597214
rect 207676 597214 207804 597216
rect 284661 597272 318932 597274
rect 284661 597216 284666 597272
rect 284722 597216 318932 597272
rect 284661 597214 318932 597216
rect 207676 597212 207723 597214
rect 207657 597211 207723 597212
rect 284661 597211 284727 597214
rect 318926 597212 318932 597214
rect 318996 597274 319002 597276
rect 428958 597274 428964 597276
rect 318996 597214 428964 597274
rect 318996 597212 319002 597214
rect 428958 597212 428964 597214
rect 429028 597212 429034 597276
rect 433333 597274 433380 597276
rect 433288 597272 433380 597274
rect 433288 597216 433338 597272
rect 433288 597214 433380 597216
rect 433333 597212 433380 597214
rect 433444 597212 433450 597276
rect 449893 597274 449959 597277
rect 450486 597274 450492 597276
rect 449893 597272 450492 597274
rect 449893 597216 449898 597272
rect 449954 597216 450492 597272
rect 449893 597214 450492 597216
rect 433333 597211 433399 597212
rect 449893 597211 449959 597214
rect 450486 597212 450492 597214
rect 450556 597212 450562 597276
rect 94037 597138 94103 597141
rect 94262 597138 94268 597140
rect 94037 597136 94268 597138
rect 94037 597080 94042 597136
rect 94098 597080 94268 597136
rect 94037 597078 94268 597080
rect 94037 597075 94103 597078
rect 94262 597076 94268 597078
rect 94332 597076 94338 597140
rect 103278 597076 103284 597140
rect 103348 597138 103354 597140
rect 103421 597138 103487 597141
rect 103348 597136 103487 597138
rect 103348 597080 103426 597136
rect 103482 597080 103487 597136
rect 103348 597078 103487 597080
rect 103348 597076 103354 597078
rect 103421 597075 103487 597078
rect 105670 597076 105676 597140
rect 105740 597138 105746 597140
rect 106181 597138 106247 597141
rect 105740 597136 106247 597138
rect 105740 597080 106186 597136
rect 106242 597080 106247 597136
rect 105740 597078 106247 597080
rect 105740 597076 105746 597078
rect 106181 597075 106247 597078
rect 106406 597076 106412 597140
rect 106476 597138 106482 597140
rect 215334 597138 215340 597140
rect 106476 597078 215340 597138
rect 106476 597076 106482 597078
rect 215334 597076 215340 597078
rect 215404 597138 215410 597140
rect 284753 597138 284819 597141
rect 434713 597140 434779 597141
rect 317638 597138 317644 597140
rect 215404 597078 219450 597138
rect 215404 597076 215410 597078
rect 99966 596940 99972 597004
rect 100036 597002 100042 597004
rect 100661 597002 100727 597005
rect 100036 597000 100727 597002
rect 100036 596944 100666 597000
rect 100722 596944 100727 597000
rect 100036 596942 100727 596944
rect 100036 596940 100042 596942
rect 100661 596939 100727 596942
rect 101070 596940 101076 597004
rect 101140 597002 101146 597004
rect 211102 597002 211108 597004
rect 101140 596942 211108 597002
rect 101140 596940 101146 596942
rect 211102 596940 211108 596942
rect 211172 597002 211178 597004
rect 212441 597002 212507 597005
rect 211172 597000 212507 597002
rect 211172 596944 212446 597000
rect 212502 596944 212507 597000
rect 211172 596942 212507 596944
rect 211172 596940 211178 596942
rect 212441 596939 212507 596942
rect 104801 596868 104867 596869
rect 104750 596804 104756 596868
rect 104820 596866 104867 596868
rect 219390 596866 219450 597078
rect 284753 597136 317644 597138
rect 284753 597080 284758 597136
rect 284814 597080 317644 597136
rect 284753 597078 317644 597080
rect 284753 597075 284819 597078
rect 317638 597076 317644 597078
rect 317708 597138 317714 597140
rect 427670 597138 427676 597140
rect 317708 597078 427676 597138
rect 317708 597076 317714 597078
rect 427670 597076 427676 597078
rect 427740 597076 427746 597140
rect 434662 597076 434668 597140
rect 434732 597138 434779 597140
rect 434732 597136 434824 597138
rect 434774 597080 434824 597136
rect 434732 597078 434824 597080
rect 434732 597076 434779 597078
rect 434713 597075 434779 597076
rect 284385 597002 284451 597005
rect 321134 597002 321140 597004
rect 284385 597000 321140 597002
rect 284385 596944 284390 597000
rect 284446 596944 321140 597000
rect 284385 596942 321140 596944
rect 284385 596939 284451 596942
rect 321134 596940 321140 596942
rect 321204 596940 321210 597004
rect 435214 597002 435220 597004
rect 325650 596942 435220 597002
rect 281809 596866 281875 596869
rect 325366 596866 325372 596868
rect 104820 596864 104912 596866
rect 104862 596808 104912 596864
rect 104820 596806 104912 596808
rect 219390 596864 325372 596866
rect 219390 596808 281814 596864
rect 281870 596808 325372 596864
rect 219390 596806 325372 596808
rect 104820 596804 104867 596806
rect 104801 596803 104867 596804
rect 281809 596803 281875 596806
rect 325366 596804 325372 596806
rect 325436 596866 325442 596868
rect 325650 596866 325710 596942
rect 435214 596940 435220 596942
rect 435284 596940 435290 597004
rect 470358 596940 470364 597004
rect 470428 597002 470434 597004
rect 470593 597002 470659 597005
rect 470428 597000 470659 597002
rect 470428 596944 470598 597000
rect 470654 596944 470659 597000
rect 470428 596942 470659 596944
rect 470428 596940 470434 596942
rect 470593 596939 470659 596942
rect 325436 596806 325710 596866
rect 325436 596804 325442 596806
rect 431718 596804 431724 596868
rect 431788 596866 431794 596868
rect 431953 596866 432019 596869
rect 431788 596864 432019 596866
rect 431788 596808 431958 596864
rect 432014 596808 432019 596864
rect 431788 596806 432019 596808
rect 431788 596804 431794 596806
rect 431953 596803 432019 596806
rect 204345 596594 204411 596597
rect 205398 596594 205404 596596
rect 204345 596592 205404 596594
rect 204345 596536 204350 596592
rect 204406 596536 205404 596592
rect 204345 596534 205404 596536
rect 204345 596531 204411 596534
rect 205398 596532 205404 596534
rect 205468 596532 205474 596596
rect 202873 596460 202939 596461
rect 202822 596396 202828 596460
rect 202892 596458 202939 596460
rect 422569 596458 422635 596461
rect 422886 596458 422892 596460
rect 202892 596456 202984 596458
rect 202934 596400 202984 596456
rect 202892 596398 202984 596400
rect 422569 596456 422892 596458
rect 422569 596400 422574 596456
rect 422630 596400 422892 596456
rect 422569 596398 422892 596400
rect 202892 596396 202939 596398
rect 202873 596395 202939 596396
rect 422569 596395 422635 596398
rect 422886 596396 422892 596398
rect 422956 596396 422962 596460
rect 95233 596322 95299 596325
rect 204253 596324 204319 596325
rect 95366 596322 95372 596324
rect 95233 596320 95372 596322
rect 95233 596264 95238 596320
rect 95294 596264 95372 596320
rect 95233 596262 95372 596264
rect 95233 596259 95299 596262
rect 95366 596260 95372 596262
rect 95436 596260 95442 596324
rect 204253 596322 204300 596324
rect 204208 596320 204300 596322
rect 204208 596264 204258 596320
rect 204208 596262 204300 596264
rect 204253 596260 204300 596262
rect 204364 596260 204370 596324
rect 311893 596322 311959 596325
rect 312854 596322 312860 596324
rect 311893 596320 312860 596322
rect 311893 596264 311898 596320
rect 311954 596264 312860 596320
rect 311893 596262 312860 596264
rect 204253 596259 204319 596260
rect 311893 596259 311959 596262
rect 312854 596260 312860 596262
rect 312924 596260 312930 596324
rect 313273 596322 313339 596325
rect 314326 596322 314332 596324
rect 313273 596320 314332 596322
rect 313273 596264 313278 596320
rect 313334 596264 314332 596320
rect 313273 596262 314332 596264
rect 313273 596259 313339 596262
rect 314326 596260 314332 596262
rect 314396 596260 314402 596324
rect 423673 596322 423739 596325
rect 424174 596322 424180 596324
rect 423673 596320 424180 596322
rect 423673 596264 423678 596320
rect 423734 596264 424180 596320
rect 423673 596262 424180 596264
rect 423673 596259 423739 596262
rect 424174 596260 424180 596262
rect 424244 596260 424250 596324
rect 425053 596322 425119 596325
rect 425278 596322 425284 596324
rect 425053 596320 425284 596322
rect 425053 596264 425058 596320
rect 425114 596264 425284 596320
rect 425053 596262 425284 596264
rect 425053 596259 425119 596262
rect 425278 596260 425284 596262
rect 425348 596260 425354 596324
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 186865 527098 186931 527101
rect 297725 527098 297791 527101
rect 407481 527098 407547 527101
rect 186865 527096 189458 527098
rect 186865 527040 186870 527096
rect 186926 527060 189458 527096
rect 297725 527096 299490 527098
rect 186926 527040 190072 527060
rect 186865 527038 190072 527040
rect 186865 527035 186931 527038
rect 78489 526690 78555 526693
rect 80002 526690 80062 527030
rect 189398 527000 190072 527038
rect 297725 527040 297730 527096
rect 297786 527060 299490 527096
rect 407481 527096 410062 527098
rect 297786 527040 300012 527060
rect 297725 527038 300012 527040
rect 297725 527035 297791 527038
rect 299430 527000 300012 527038
rect 407481 527040 407486 527096
rect 407542 527040 410062 527096
rect 407481 527038 410062 527040
rect 407481 527035 407547 527038
rect 410002 527030 410062 527038
rect 78489 526688 80062 526690
rect 78489 526632 78494 526688
rect 78550 526632 80062 526688
rect 78489 526630 80062 526632
rect 78489 526627 78555 526630
rect 78305 526554 78371 526557
rect 407665 526554 407731 526557
rect 78305 526552 80062 526554
rect 78305 526496 78310 526552
rect 78366 526496 80062 526552
rect 78305 526494 80062 526496
rect 78305 526491 78371 526494
rect 80002 525942 80062 526494
rect 407665 526552 410062 526554
rect 407665 526496 407670 526552
rect 407726 526496 410062 526552
rect 407665 526494 410062 526496
rect 407665 526491 407731 526494
rect 186681 526010 186747 526013
rect 189073 526010 189139 526013
rect 298001 526010 298067 526013
rect 186681 526008 189458 526010
rect 186681 525952 186686 526008
rect 186742 525952 189078 526008
rect 189134 525972 189458 526008
rect 298001 526008 299490 526010
rect 189134 525952 190072 525972
rect 186681 525950 190072 525952
rect 186681 525947 186747 525950
rect 189073 525947 189139 525950
rect 189398 525912 190072 525950
rect 298001 525952 298006 526008
rect 298062 525972 299490 526008
rect 298062 525952 300012 525972
rect 298001 525950 300012 525952
rect 298001 525947 298067 525950
rect 299430 525912 300012 525950
rect 410002 525942 410062 526494
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 187325 524378 187391 524381
rect 188337 524378 188403 524381
rect 298001 524378 298067 524381
rect 187325 524376 189458 524378
rect 187325 524320 187330 524376
rect 187386 524320 188342 524376
rect 188398 524340 189458 524376
rect 298001 524376 299490 524378
rect 188398 524320 190072 524340
rect 187325 524318 190072 524320
rect 187325 524315 187391 524318
rect 188337 524315 188403 524318
rect 78305 523698 78371 523701
rect 80002 523698 80062 524310
rect 189398 524280 190072 524318
rect 298001 524320 298006 524376
rect 298062 524340 299490 524376
rect 583520 524364 584960 524454
rect 298062 524320 300012 524340
rect 298001 524318 300012 524320
rect 298001 524315 298067 524318
rect 299430 524280 300012 524318
rect 78305 523696 80062 523698
rect 78305 523640 78310 523696
rect 78366 523640 80062 523696
rect 78305 523638 80062 523640
rect 78305 523635 78371 523638
rect 407798 523636 407804 523700
rect 407868 523698 407874 523700
rect 410002 523698 410062 524310
rect 407868 523638 410062 523698
rect 407868 523636 407874 523638
rect 77569 523290 77635 523293
rect 77937 523290 78003 523293
rect 187417 523290 187483 523293
rect 187785 523290 187851 523293
rect 297909 523290 297975 523293
rect 407665 523290 407731 523293
rect 408033 523290 408099 523293
rect 77569 523288 80062 523290
rect 77569 523232 77574 523288
rect 77630 523232 77942 523288
rect 77998 523232 80062 523288
rect 77569 523230 80062 523232
rect 77569 523227 77635 523230
rect 77937 523227 78003 523230
rect 80002 523222 80062 523230
rect 187417 523288 189458 523290
rect 187417 523232 187422 523288
rect 187478 523232 187790 523288
rect 187846 523252 189458 523288
rect 297909 523288 299490 523290
rect 187846 523232 190072 523252
rect 187417 523230 190072 523232
rect 187417 523227 187483 523230
rect 187785 523227 187851 523230
rect 189398 523192 190072 523230
rect 297909 523232 297914 523288
rect 297970 523252 299490 523288
rect 407665 523288 410062 523290
rect 297970 523232 300012 523252
rect 297909 523230 300012 523232
rect 297909 523227 297975 523230
rect 299430 523192 300012 523230
rect 407665 523232 407670 523288
rect 407726 523232 408038 523288
rect 408094 523232 410062 523288
rect 407665 523230 410062 523232
rect 407665 523227 407731 523230
rect 408033 523227 408099 523230
rect 410002 523222 410062 523230
rect 187233 521658 187299 521661
rect 187969 521658 188035 521661
rect 297449 521658 297515 521661
rect 187233 521656 189458 521658
rect 187233 521600 187238 521656
rect 187294 521600 187974 521656
rect 188030 521620 189458 521656
rect 297449 521656 299490 521658
rect 188030 521600 190072 521620
rect 187233 521598 190072 521600
rect 187233 521595 187299 521598
rect 187969 521595 188035 521598
rect 78121 520978 78187 520981
rect 80002 520978 80062 521590
rect 189398 521560 190072 521598
rect 297449 521600 297454 521656
rect 297510 521620 299490 521656
rect 297510 521600 300012 521620
rect 297449 521598 300012 521600
rect 297449 521595 297515 521598
rect 299430 521560 300012 521598
rect 78121 520976 80062 520978
rect 78121 520920 78126 520976
rect 78182 520920 80062 520976
rect 78121 520918 80062 520920
rect 407573 520978 407639 520981
rect 410002 520978 410062 521590
rect 407573 520976 410062 520978
rect 407573 520920 407578 520976
rect 407634 520920 410062 520976
rect 407573 520918 410062 520920
rect 78121 520915 78187 520918
rect 407573 520915 407639 520918
rect 77753 520298 77819 520301
rect 188153 520298 188219 520301
rect 297817 520298 297883 520301
rect 408125 520298 408191 520301
rect 77753 520296 80062 520298
rect 77753 520240 77758 520296
rect 77814 520240 80062 520296
rect 77753 520238 80062 520240
rect 77753 520235 77819 520238
rect 80002 520230 80062 520238
rect 188153 520296 190010 520298
rect 188153 520240 188158 520296
rect 188214 520260 190010 520296
rect 297817 520296 299858 520298
rect 188214 520240 190072 520260
rect 188153 520238 190072 520240
rect 188153 520235 188219 520238
rect 189950 520200 190072 520238
rect 297817 520240 297822 520296
rect 297878 520260 299858 520296
rect 408125 520296 410062 520298
rect 297878 520240 300012 520260
rect 297817 520238 300012 520240
rect 297817 520235 297883 520238
rect 299798 520200 300012 520238
rect 408125 520240 408130 520296
rect 408186 520240 410062 520296
rect 408125 520238 410062 520240
rect 408125 520235 408191 520238
rect 410002 520230 410062 520238
rect 188061 518666 188127 518669
rect 297541 518666 297607 518669
rect 188061 518664 189458 518666
rect 188061 518608 188066 518664
rect 188122 518628 189458 518664
rect 297541 518664 299490 518666
rect 188122 518608 190072 518628
rect 188061 518606 190072 518608
rect 188061 518603 188127 518606
rect 78029 517986 78095 517989
rect 80002 517986 80062 518598
rect 189398 518568 190072 518606
rect 297541 518608 297546 518664
rect 297602 518628 299490 518664
rect 297602 518608 300012 518628
rect 297541 518606 300012 518608
rect 297541 518603 297607 518606
rect 299430 518568 300012 518606
rect 78029 517984 80062 517986
rect 78029 517928 78034 517984
rect 78090 517928 80062 517984
rect 78029 517926 80062 517928
rect 407481 517986 407547 517989
rect 410002 517986 410062 518598
rect 407481 517984 410062 517986
rect 407481 517928 407486 517984
rect 407542 517928 410062 517984
rect 407481 517926 410062 517928
rect 78029 517923 78095 517926
rect 407481 517923 407547 517926
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 296989 500850 297055 500853
rect 297909 500850 297975 500853
rect 296989 500848 297975 500850
rect 296989 500792 296994 500848
rect 297050 500792 297914 500848
rect 297970 500792 297975 500848
rect 296989 500790 297975 500792
rect 296989 500787 297055 500790
rect 297909 500787 297975 500790
rect 187049 500306 187115 500309
rect 297909 500306 297975 500309
rect 408401 500306 408467 500309
rect 187049 500304 189458 500306
rect 187049 500248 187054 500304
rect 187110 500268 189458 500304
rect 297909 500304 299490 500306
rect 187110 500248 190072 500268
rect 187049 500246 190072 500248
rect 187049 500243 187115 500246
rect 78581 499898 78647 499901
rect 80002 499898 80062 500238
rect 189398 500208 190072 500246
rect 297909 500248 297914 500304
rect 297970 500268 299490 500304
rect 408401 500304 410062 500306
rect 297970 500248 300012 500268
rect 297909 500246 300012 500248
rect 297909 500243 297975 500246
rect 299430 500208 300012 500246
rect 408401 500248 408406 500304
rect 408462 500248 410062 500304
rect 408401 500246 410062 500248
rect 408401 500243 408467 500246
rect 410002 500238 410062 500246
rect 78581 499896 80062 499898
rect 78581 499840 78586 499896
rect 78642 499840 80062 499896
rect 78581 499838 80062 499840
rect 78581 499835 78647 499838
rect 77937 498674 78003 498677
rect 187601 498674 187667 498677
rect 297449 498674 297515 498677
rect 408309 498674 408375 498677
rect 77937 498672 80062 498674
rect 77937 498616 77942 498672
rect 77998 498616 80062 498672
rect 77937 498614 80062 498616
rect 77937 498611 78003 498614
rect 80002 498606 80062 498614
rect 187601 498672 189458 498674
rect 187601 498616 187606 498672
rect 187662 498636 189458 498672
rect 297449 498672 299490 498674
rect 187662 498616 190072 498636
rect 187601 498614 190072 498616
rect 187601 498611 187667 498614
rect 189398 498576 190072 498614
rect 297449 498616 297454 498672
rect 297510 498636 299490 498672
rect 408309 498672 410062 498674
rect 297510 498616 300012 498636
rect 297449 498614 300012 498616
rect 297449 498611 297515 498614
rect 299430 498576 300012 498614
rect 408309 498616 408314 498672
rect 408370 498616 410062 498672
rect 408309 498614 410062 498616
rect 408309 498611 408375 498614
rect 410002 498606 410062 498614
rect 77661 498402 77727 498405
rect 407849 498402 407915 498405
rect 77661 498400 79426 498402
rect 77661 498344 77666 498400
rect 77722 498364 79426 498400
rect 407849 498400 409522 498402
rect 77722 498344 80032 498364
rect 77661 498342 80032 498344
rect 77661 498339 77727 498342
rect 79366 498304 80032 498342
rect 189398 498304 190072 498364
rect 299430 498304 300012 498364
rect 407849 498344 407854 498400
rect 407910 498364 409522 498400
rect 407910 498344 410032 498364
rect 407849 498342 410032 498344
rect 407849 498339 407915 498342
rect 409462 498304 410032 498342
rect 186589 498266 186655 498269
rect 187049 498266 187115 498269
rect 189398 498266 189458 498304
rect 186589 498264 189458 498266
rect 186589 498208 186594 498264
rect 186650 498208 187054 498264
rect 187110 498208 189458 498264
rect 186589 498206 189458 498208
rect 296897 498266 296963 498269
rect 297817 498266 297883 498269
rect 299430 498266 299490 498304
rect 296897 498264 299490 498266
rect 296897 498208 296902 498264
rect 296958 498208 297822 498264
rect 297878 498208 299490 498264
rect 296897 498206 299490 498208
rect 408033 498266 408099 498269
rect 408309 498266 408375 498269
rect 408033 498264 408375 498266
rect 408033 498208 408038 498264
rect 408094 498208 408314 498264
rect 408370 498208 408375 498264
rect 408033 498206 408375 498208
rect 186589 498203 186655 498206
rect 187049 498203 187115 498206
rect 296897 498203 296963 498206
rect 297817 498203 297883 498206
rect 408033 498203 408099 498206
rect 408309 498203 408375 498206
rect 583520 497844 584960 498084
rect 285581 489834 285647 489837
rect 407798 489834 407804 489836
rect 285581 489832 407804 489834
rect 285581 489776 285586 489832
rect 285642 489776 407804 489832
rect 285581 489774 407804 489776
rect 285581 489771 285647 489774
rect 407798 489772 407804 489774
rect 407868 489772 407874 489836
rect 110505 489428 110571 489429
rect 110454 489426 110460 489428
rect 110414 489366 110460 489426
rect 110524 489424 110571 489428
rect 110566 489368 110571 489424
rect 110454 489364 110460 489366
rect 110524 489364 110571 489368
rect 110505 489363 110571 489364
rect 325325 489156 325391 489157
rect 325325 489152 325372 489156
rect 325436 489154 325442 489156
rect 325325 489096 325330 489152
rect 325325 489092 325372 489096
rect 325436 489094 325482 489154
rect 325436 489092 325442 489094
rect 325325 489091 325391 489092
rect -960 488596 480 488836
rect 285029 488610 285095 488613
rect 285581 488610 285647 488613
rect 285029 488608 285647 488610
rect 285029 488552 285034 488608
rect 285090 488552 285586 488608
rect 285642 488552 285647 488608
rect 285029 488550 285647 488552
rect 285029 488547 285095 488550
rect 285581 488547 285647 488550
rect 92933 488476 92999 488477
rect 94221 488476 94287 488477
rect 97809 488476 97875 488477
rect 92933 488472 92980 488476
rect 93044 488474 93050 488476
rect 92933 488416 92938 488472
rect 92933 488412 92980 488416
rect 93044 488414 93090 488474
rect 94221 488472 94268 488476
rect 94332 488474 94338 488476
rect 97758 488474 97764 488476
rect 94221 488416 94226 488472
rect 93044 488412 93050 488414
rect 94221 488412 94268 488416
rect 94332 488414 94378 488474
rect 97718 488414 97764 488474
rect 97828 488472 97875 488476
rect 97870 488416 97875 488472
rect 94332 488412 94338 488414
rect 97758 488412 97764 488414
rect 97828 488412 97875 488416
rect 98862 488412 98868 488476
rect 98932 488474 98938 488476
rect 99189 488474 99255 488477
rect 100017 488476 100083 488477
rect 101121 488476 101187 488477
rect 102409 488476 102475 488477
rect 104801 488476 104867 488477
rect 105353 488476 105419 488477
rect 105721 488476 105787 488477
rect 115657 488476 115723 488477
rect 120625 488476 120691 488477
rect 125593 488476 125659 488477
rect 99966 488474 99972 488476
rect 98932 488472 99255 488474
rect 98932 488416 99194 488472
rect 99250 488416 99255 488472
rect 98932 488414 99255 488416
rect 99926 488414 99972 488474
rect 100036 488472 100083 488476
rect 101070 488474 101076 488476
rect 100078 488416 100083 488472
rect 98932 488412 98938 488414
rect 92933 488411 92999 488412
rect 94221 488411 94287 488412
rect 97809 488411 97875 488412
rect 99189 488411 99255 488414
rect 99966 488412 99972 488414
rect 100036 488412 100083 488416
rect 101030 488414 101076 488474
rect 101140 488472 101187 488476
rect 102358 488474 102364 488476
rect 101182 488416 101187 488472
rect 101070 488412 101076 488414
rect 101140 488412 101187 488416
rect 102318 488414 102364 488474
rect 102428 488472 102475 488476
rect 104750 488474 104756 488476
rect 102470 488416 102475 488472
rect 102358 488412 102364 488414
rect 102428 488412 102475 488416
rect 104710 488414 104756 488474
rect 104820 488472 104867 488476
rect 105302 488474 105308 488476
rect 104862 488416 104867 488472
rect 104750 488412 104756 488414
rect 104820 488412 104867 488416
rect 105262 488414 105308 488474
rect 105372 488472 105419 488476
rect 105670 488474 105676 488476
rect 105414 488416 105419 488472
rect 105302 488412 105308 488414
rect 105372 488412 105419 488416
rect 105630 488414 105676 488474
rect 105740 488472 105787 488476
rect 115606 488474 115612 488476
rect 105782 488416 105787 488472
rect 105670 488412 105676 488414
rect 105740 488412 105787 488416
rect 115566 488414 115612 488474
rect 115676 488472 115723 488476
rect 120574 488474 120580 488476
rect 115718 488416 115723 488472
rect 115606 488412 115612 488414
rect 115676 488412 115723 488416
rect 120534 488414 120580 488474
rect 120644 488472 120691 488476
rect 125542 488474 125548 488476
rect 120686 488416 120691 488472
rect 120574 488412 120580 488414
rect 120644 488412 120691 488416
rect 125502 488414 125548 488474
rect 125612 488472 125659 488476
rect 125654 488416 125659 488472
rect 125542 488412 125548 488414
rect 125612 488412 125659 488416
rect 130510 488412 130516 488476
rect 130580 488474 130586 488476
rect 130653 488474 130719 488477
rect 135529 488476 135595 488477
rect 140681 488476 140747 488477
rect 215293 488476 215359 488477
rect 135478 488474 135484 488476
rect 130580 488472 130719 488474
rect 130580 488416 130658 488472
rect 130714 488416 130719 488472
rect 130580 488414 130719 488416
rect 135438 488414 135484 488474
rect 135548 488472 135595 488476
rect 140630 488474 140636 488476
rect 135590 488416 135595 488472
rect 130580 488412 130586 488414
rect 100017 488411 100083 488412
rect 101121 488411 101187 488412
rect 102409 488411 102475 488412
rect 104801 488411 104867 488412
rect 105353 488411 105419 488412
rect 105721 488411 105787 488412
rect 115657 488411 115723 488412
rect 120625 488411 120691 488412
rect 125593 488411 125659 488412
rect 130653 488411 130719 488414
rect 135478 488412 135484 488414
rect 135548 488412 135595 488416
rect 140590 488414 140636 488474
rect 140700 488472 140747 488476
rect 205398 488474 205404 488476
rect 140742 488416 140747 488472
rect 140630 488412 140636 488414
rect 140700 488412 140747 488416
rect 135529 488411 135595 488412
rect 140681 488411 140747 488412
rect 190410 488414 205404 488474
rect 95325 488340 95391 488341
rect 95325 488338 95372 488340
rect 95244 488336 95372 488338
rect 95436 488338 95442 488340
rect 188889 488338 188955 488341
rect 190410 488338 190470 488414
rect 205398 488412 205404 488414
rect 205468 488412 205474 488476
rect 215293 488472 215340 488476
rect 215404 488474 215410 488476
rect 215293 488416 215298 488472
rect 215293 488412 215340 488416
rect 215404 488414 215450 488474
rect 215404 488412 215410 488414
rect 220486 488412 220492 488476
rect 220556 488474 220562 488476
rect 220721 488474 220787 488477
rect 220556 488472 220787 488474
rect 220556 488416 220726 488472
rect 220782 488416 220787 488472
rect 220556 488414 220787 488416
rect 220556 488412 220562 488414
rect 215293 488411 215359 488412
rect 220721 488411 220787 488414
rect 225454 488412 225460 488476
rect 225524 488474 225530 488476
rect 226241 488474 226307 488477
rect 230473 488476 230539 488477
rect 230422 488474 230428 488476
rect 225524 488472 226307 488474
rect 225524 488416 226246 488472
rect 226302 488416 226307 488472
rect 225524 488414 226307 488416
rect 230382 488414 230428 488474
rect 230492 488472 230539 488476
rect 230534 488416 230539 488472
rect 225524 488412 225530 488414
rect 226241 488411 226307 488414
rect 230422 488412 230428 488414
rect 230492 488412 230539 488416
rect 230473 488411 230539 488412
rect 330477 488476 330543 488477
rect 335445 488476 335511 488477
rect 340597 488476 340663 488477
rect 330477 488472 330524 488476
rect 330588 488474 330594 488476
rect 330477 488416 330482 488472
rect 330477 488412 330524 488416
rect 330588 488414 330634 488474
rect 335445 488472 335492 488476
rect 335556 488474 335562 488476
rect 335445 488416 335450 488472
rect 330588 488412 330594 488414
rect 335445 488412 335492 488416
rect 335556 488414 335602 488474
rect 340597 488472 340644 488476
rect 340708 488474 340714 488476
rect 340597 488416 340602 488472
rect 335556 488412 335562 488414
rect 340597 488412 340644 488416
rect 340708 488414 340754 488474
rect 340708 488412 340714 488414
rect 345606 488412 345612 488476
rect 345676 488474 345682 488476
rect 345749 488474 345815 488477
rect 345676 488472 345815 488474
rect 345676 488416 345754 488472
rect 345810 488416 345815 488472
rect 345676 488414 345815 488416
rect 345676 488412 345682 488414
rect 330477 488411 330543 488412
rect 335445 488411 335511 488412
rect 340597 488411 340663 488412
rect 345749 488411 345815 488414
rect 350349 488476 350415 488477
rect 350349 488472 350396 488476
rect 350460 488474 350466 488476
rect 350349 488416 350354 488472
rect 350349 488412 350396 488416
rect 350460 488414 350506 488474
rect 350460 488412 350466 488414
rect 355542 488412 355548 488476
rect 355612 488474 355618 488476
rect 355777 488474 355843 488477
rect 355612 488472 355843 488474
rect 355612 488416 355782 488472
rect 355838 488416 355843 488472
rect 355612 488414 355843 488416
rect 355612 488412 355618 488414
rect 350349 488411 350415 488412
rect 355777 488411 355843 488414
rect 360469 488476 360535 488477
rect 360469 488472 360516 488476
rect 360580 488474 360586 488476
rect 422569 488474 422635 488477
rect 422886 488474 422892 488476
rect 360469 488416 360474 488472
rect 360469 488412 360516 488416
rect 360580 488414 360626 488474
rect 422569 488472 422892 488474
rect 422569 488416 422574 488472
rect 422630 488416 422892 488472
rect 422569 488414 422892 488416
rect 360580 488412 360586 488414
rect 360469 488411 360535 488412
rect 422569 488411 422635 488414
rect 422886 488412 422892 488414
rect 422956 488412 422962 488476
rect 423673 488474 423739 488477
rect 424174 488474 424180 488476
rect 423673 488472 424180 488474
rect 423673 488416 423678 488472
rect 423734 488416 424180 488472
rect 423673 488414 424180 488416
rect 423673 488411 423739 488414
rect 424174 488412 424180 488414
rect 424244 488412 424250 488476
rect 434713 488474 434779 488477
rect 435214 488474 435220 488476
rect 434713 488472 435220 488474
rect 434713 488416 434718 488472
rect 434774 488416 435220 488472
rect 434713 488414 435220 488416
rect 434713 488411 434779 488414
rect 435214 488412 435220 488414
rect 435284 488412 435290 488476
rect 440233 488474 440299 488477
rect 440366 488474 440372 488476
rect 440233 488472 440372 488474
rect 440233 488416 440238 488472
rect 440294 488416 440372 488472
rect 440233 488414 440372 488416
rect 440233 488411 440299 488414
rect 440366 488412 440372 488414
rect 440436 488412 440442 488476
rect 444373 488474 444439 488477
rect 445518 488474 445524 488476
rect 444373 488472 445524 488474
rect 444373 488416 444378 488472
rect 444434 488416 445524 488472
rect 444373 488414 445524 488416
rect 444373 488411 444439 488414
rect 445518 488412 445524 488414
rect 445588 488412 445594 488476
rect 449893 488474 449959 488477
rect 450486 488474 450492 488476
rect 449893 488472 450492 488474
rect 449893 488416 449898 488472
rect 449954 488416 450492 488472
rect 449893 488414 450492 488416
rect 449893 488411 449959 488414
rect 450486 488412 450492 488414
rect 450556 488412 450562 488476
rect 95436 488336 190470 488338
rect 95244 488280 95330 488336
rect 95436 488280 188894 488336
rect 188950 488280 190470 488336
rect 95244 488278 95372 488280
rect 95325 488276 95372 488278
rect 95436 488278 190470 488280
rect 313917 488338 313983 488341
rect 314326 488338 314332 488340
rect 313917 488336 314332 488338
rect 313917 488280 313922 488336
rect 313978 488280 314332 488336
rect 313917 488278 314332 488280
rect 95436 488276 95442 488278
rect 95325 488275 95391 488276
rect 188889 488275 188955 488278
rect 313917 488275 313983 488278
rect 314326 488276 314332 488278
rect 314396 488338 314402 488340
rect 407941 488338 408007 488341
rect 425278 488338 425284 488340
rect 314396 488336 408007 488338
rect 314396 488280 407946 488336
rect 408002 488280 408007 488336
rect 314396 488278 408007 488280
rect 314396 488276 314402 488278
rect 407941 488275 408007 488278
rect 412590 488278 425284 488338
rect 315297 488202 315363 488205
rect 315430 488202 315436 488204
rect 315297 488200 315436 488202
rect 315297 488144 315302 488200
rect 315358 488144 315436 488200
rect 315297 488142 315436 488144
rect 315297 488139 315363 488142
rect 315430 488140 315436 488142
rect 315500 488202 315506 488204
rect 407757 488202 407823 488205
rect 412590 488202 412650 488278
rect 425278 488276 425284 488278
rect 425348 488276 425354 488340
rect 430573 488338 430639 488341
rect 430982 488338 430988 488340
rect 430573 488336 430988 488338
rect 430573 488280 430578 488336
rect 430634 488280 430988 488336
rect 430573 488278 430988 488280
rect 430573 488275 430639 488278
rect 430982 488276 430988 488278
rect 431052 488276 431058 488340
rect 465073 488338 465139 488341
rect 465390 488338 465396 488340
rect 465073 488336 465396 488338
rect 465073 488280 465078 488336
rect 465134 488280 465396 488336
rect 465073 488278 465396 488280
rect 465073 488275 465139 488278
rect 465390 488276 465396 488278
rect 465460 488276 465466 488340
rect 315500 488200 412650 488202
rect 315500 488144 407762 488200
rect 407818 488144 412650 488200
rect 315500 488142 412650 488144
rect 427813 488202 427879 488205
rect 428958 488202 428964 488204
rect 427813 488200 428964 488202
rect 427813 488144 427818 488200
rect 427874 488144 428964 488200
rect 427813 488142 428964 488144
rect 315500 488140 315506 488142
rect 407757 488139 407823 488142
rect 427813 488139 427879 488142
rect 428958 488140 428964 488142
rect 429028 488140 429034 488204
rect 429193 488202 429259 488205
rect 429878 488202 429884 488204
rect 429193 488200 429884 488202
rect 429193 488144 429198 488200
rect 429254 488144 429884 488200
rect 429193 488142 429884 488144
rect 429193 488139 429259 488142
rect 429878 488140 429884 488142
rect 429948 488140 429954 488204
rect 434713 488202 434779 488205
rect 435582 488202 435588 488204
rect 434713 488200 435588 488202
rect 434713 488144 434718 488200
rect 434774 488144 435588 488200
rect 434713 488142 435588 488144
rect 434713 488139 434779 488142
rect 435582 488140 435588 488142
rect 435652 488140 435658 488204
rect 202873 488066 202939 488069
rect 204253 488068 204319 488069
rect 203006 488066 203012 488068
rect 202873 488064 203012 488066
rect 202873 488008 202878 488064
rect 202934 488008 203012 488064
rect 202873 488006 203012 488008
rect 202873 488003 202939 488006
rect 203006 488004 203012 488006
rect 203076 488004 203082 488068
rect 204253 488066 204300 488068
rect 204208 488064 204300 488066
rect 204208 488008 204258 488064
rect 204208 488006 204300 488008
rect 204253 488004 204300 488006
rect 204364 488004 204370 488068
rect 211797 488066 211863 488069
rect 212206 488066 212212 488068
rect 211797 488064 212212 488066
rect 211797 488008 211802 488064
rect 211858 488008 212212 488064
rect 211797 488006 212212 488008
rect 204253 488003 204319 488004
rect 211797 488003 211863 488006
rect 212206 488004 212212 488006
rect 212276 488004 212282 488068
rect 282361 488066 282427 488069
rect 407481 488066 407547 488069
rect 455413 488068 455479 488069
rect 455413 488066 455460 488068
rect 282361 488064 407547 488066
rect 282361 488008 282366 488064
rect 282422 488008 407486 488064
rect 407542 488008 407547 488064
rect 282361 488006 407547 488008
rect 455368 488064 455460 488066
rect 455368 488008 455418 488064
rect 455368 488006 455460 488008
rect 282361 488003 282427 488006
rect 407481 488003 407547 488006
rect 455413 488004 455460 488006
rect 455524 488004 455530 488068
rect 470593 488066 470659 488069
rect 470726 488066 470732 488068
rect 470593 488064 470732 488066
rect 470593 488008 470598 488064
rect 470654 488008 470732 488064
rect 470593 488006 470732 488008
rect 455413 488003 455479 488004
rect 470593 488003 470659 488006
rect 470726 488004 470732 488006
rect 470796 488004 470802 488068
rect 211153 487932 211219 487933
rect 235625 487932 235691 487933
rect 211102 487930 211108 487932
rect 211062 487870 211108 487930
rect 211172 487928 211219 487932
rect 235574 487930 235580 487932
rect 211214 487872 211219 487928
rect 211102 487868 211108 487870
rect 211172 487868 211219 487872
rect 235534 487870 235580 487930
rect 235644 487928 235691 487932
rect 235686 487872 235691 487928
rect 235574 487868 235580 487870
rect 235644 487868 235691 487872
rect 240542 487868 240548 487932
rect 240612 487930 240618 487932
rect 241421 487930 241487 487933
rect 240612 487928 241487 487930
rect 240612 487872 241426 487928
rect 241482 487872 241487 487928
rect 240612 487870 241487 487872
rect 240612 487868 240618 487870
rect 211153 487867 211219 487868
rect 235625 487867 235691 487868
rect 241421 487867 241487 487870
rect 318885 487932 318951 487933
rect 318885 487928 318932 487932
rect 318996 487930 319002 487932
rect 459553 487930 459619 487933
rect 460422 487930 460428 487932
rect 318885 487872 318890 487928
rect 318885 487868 318932 487872
rect 318996 487870 319042 487930
rect 459553 487928 460428 487930
rect 459553 487872 459558 487928
rect 459614 487872 460428 487928
rect 459553 487870 460428 487872
rect 318996 487868 319002 487870
rect 318885 487867 318951 487868
rect 459553 487867 459619 487870
rect 460422 487868 460428 487870
rect 460492 487868 460498 487932
rect 189901 487794 189967 487797
rect 219893 487794 219959 487797
rect 189901 487792 219959 487794
rect 189901 487736 189906 487792
rect 189962 487736 219898 487792
rect 219954 487736 219959 487792
rect 189901 487734 219959 487736
rect 189901 487731 189967 487734
rect 219893 487731 219959 487734
rect 426433 487794 426499 487797
rect 427670 487794 427676 487796
rect 426433 487792 427676 487794
rect 426433 487736 426438 487792
rect 426494 487736 427676 487792
rect 426433 487734 427676 487736
rect 426433 487731 426499 487734
rect 427670 487732 427676 487734
rect 427740 487732 427746 487796
rect 432045 487658 432111 487661
rect 432270 487658 432276 487660
rect 432045 487656 432276 487658
rect 432045 487600 432050 487656
rect 432106 487600 432276 487656
rect 432045 487598 432276 487600
rect 432045 487595 432111 487598
rect 432270 487596 432276 487598
rect 432340 487596 432346 487660
rect 103278 487460 103284 487524
rect 103348 487522 103354 487524
rect 103421 487522 103487 487525
rect 210049 487524 210115 487525
rect 209998 487522 210004 487524
rect 103348 487520 103487 487522
rect 103348 487464 103426 487520
rect 103482 487464 103487 487520
rect 103348 487462 103487 487464
rect 209958 487462 210004 487522
rect 210068 487520 210115 487524
rect 210110 487464 210115 487520
rect 103348 487460 103354 487462
rect 103421 487459 103487 487462
rect 209998 487460 210004 487462
rect 210068 487460 210115 487464
rect 210049 487459 210115 487460
rect 213177 487522 213243 487525
rect 250437 487524 250503 487525
rect 213310 487522 213316 487524
rect 213177 487520 213316 487522
rect 213177 487464 213182 487520
rect 213238 487464 213316 487520
rect 213177 487462 213316 487464
rect 213177 487459 213243 487462
rect 213310 487460 213316 487462
rect 213380 487460 213386 487524
rect 250437 487520 250484 487524
rect 250548 487522 250554 487524
rect 250437 487464 250442 487520
rect 250437 487460 250484 487464
rect 250548 487462 250594 487522
rect 250548 487460 250554 487462
rect 250437 487459 250503 487460
rect 204897 487386 204963 487389
rect 245561 487388 245627 487389
rect 205398 487386 205404 487388
rect 204897 487384 205404 487386
rect 204897 487328 204902 487384
rect 204958 487328 205404 487384
rect 204897 487326 205404 487328
rect 204897 487323 204963 487326
rect 205398 487324 205404 487326
rect 205468 487324 205474 487388
rect 245510 487386 245516 487388
rect 245470 487326 245516 487386
rect 245580 487384 245627 487388
rect 245622 487328 245627 487384
rect 245510 487324 245516 487326
rect 245580 487324 245627 487328
rect 323342 487324 323348 487388
rect 323412 487386 323418 487388
rect 323577 487386 323643 487389
rect 433333 487388 433399 487389
rect 433333 487386 433380 487388
rect 323412 487384 323643 487386
rect 323412 487328 323582 487384
rect 323638 487328 323643 487384
rect 323412 487326 323643 487328
rect 433288 487384 433380 487386
rect 433288 487328 433338 487384
rect 433288 487326 433380 487328
rect 323412 487324 323418 487326
rect 245561 487323 245627 487324
rect 323577 487323 323643 487326
rect 433333 487324 433380 487326
rect 433444 487324 433450 487388
rect 433333 487323 433399 487324
rect 203006 487188 203012 487252
rect 203076 487250 203082 487252
rect 203517 487250 203583 487253
rect 203076 487248 203583 487250
rect 203076 487192 203522 487248
rect 203578 487192 203583 487248
rect 203076 487190 203583 487192
rect 203076 487188 203082 487190
rect 203517 487187 203583 487190
rect 204294 487188 204300 487252
rect 204364 487250 204370 487252
rect 205081 487250 205147 487253
rect 207657 487252 207723 487253
rect 207606 487250 207612 487252
rect 204364 487248 205147 487250
rect 204364 487192 205086 487248
rect 205142 487192 205147 487248
rect 204364 487190 205147 487192
rect 207566 487190 207612 487250
rect 207676 487248 207723 487252
rect 207718 487192 207723 487248
rect 204364 487188 204370 487190
rect 205081 487187 205147 487190
rect 207606 487188 207612 487190
rect 207676 487188 207723 487192
rect 208894 487188 208900 487252
rect 208964 487250 208970 487252
rect 209037 487250 209103 487253
rect 208964 487248 209103 487250
rect 208964 487192 209042 487248
rect 209098 487192 209103 487248
rect 208964 487190 209103 487192
rect 208964 487188 208970 487190
rect 207657 487187 207723 487188
rect 209037 487187 209103 487190
rect 214557 487250 214623 487253
rect 214782 487250 214788 487252
rect 214557 487248 214788 487250
rect 214557 487192 214562 487248
rect 214618 487192 214788 487248
rect 214557 487190 214788 487192
rect 214557 487187 214623 487190
rect 214782 487188 214788 487190
rect 214852 487188 214858 487252
rect 215702 487188 215708 487252
rect 215772 487250 215778 487252
rect 215937 487250 216003 487253
rect 215772 487248 216003 487250
rect 215772 487192 215942 487248
rect 215998 487192 216003 487248
rect 215772 487190 216003 487192
rect 215772 487188 215778 487190
rect 215937 487187 216003 487190
rect 312537 487250 312603 487253
rect 312854 487250 312860 487252
rect 312537 487248 312860 487250
rect 312537 487192 312542 487248
rect 312598 487192 312860 487248
rect 312537 487190 312860 487192
rect 312537 487187 312603 487190
rect 312854 487188 312860 487190
rect 312924 487188 312930 487252
rect 317638 487188 317644 487252
rect 317708 487250 317714 487252
rect 318057 487250 318123 487253
rect 317708 487248 318123 487250
rect 317708 487192 318062 487248
rect 318118 487192 318123 487248
rect 317708 487190 318123 487192
rect 317708 487188 317714 487190
rect 318057 487187 318123 487190
rect 319437 487250 319503 487253
rect 320081 487252 320147 487253
rect 320030 487250 320036 487252
rect 319437 487248 320036 487250
rect 320100 487250 320147 487252
rect 320817 487250 320883 487253
rect 322197 487252 322263 487253
rect 324865 487252 324931 487253
rect 321134 487250 321140 487252
rect 320100 487248 320228 487250
rect 319437 487192 319442 487248
rect 319498 487192 320036 487248
rect 320142 487192 320228 487248
rect 319437 487190 320036 487192
rect 319437 487187 319503 487190
rect 320030 487188 320036 487190
rect 320100 487190 320228 487192
rect 320817 487248 321140 487250
rect 320817 487192 320822 487248
rect 320878 487192 321140 487248
rect 320817 487190 321140 487192
rect 320100 487188 320147 487190
rect 320081 487187 320147 487188
rect 320817 487187 320883 487190
rect 321134 487188 321140 487190
rect 321204 487188 321210 487252
rect 322197 487248 322244 487252
rect 322308 487250 322314 487252
rect 324814 487250 324820 487252
rect 322197 487192 322202 487248
rect 322197 487188 322244 487192
rect 322308 487190 322354 487250
rect 324774 487190 324820 487250
rect 324884 487248 324931 487252
rect 324926 487192 324931 487248
rect 322308 487188 322314 487190
rect 324814 487188 324820 487190
rect 324884 487188 324931 487192
rect 325734 487188 325740 487252
rect 325804 487250 325810 487252
rect 326337 487250 326403 487253
rect 325804 487248 326403 487250
rect 325804 487192 326342 487248
rect 326398 487192 326403 487248
rect 325804 487190 326403 487192
rect 325804 487188 325810 487190
rect 322197 487187 322263 487188
rect 324865 487187 324931 487188
rect 326337 487187 326403 487190
rect 434713 487250 434779 487253
rect 434846 487250 434852 487252
rect 434713 487248 434852 487250
rect 434713 487192 434718 487248
rect 434774 487192 434852 487248
rect 434713 487190 434852 487192
rect 434713 487187 434779 487190
rect 434846 487188 434852 487190
rect 434916 487188 434922 487252
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 219709 476778 219775 476781
rect 282126 476778 282132 476780
rect 219709 476776 282132 476778
rect 219709 476720 219714 476776
rect 219770 476720 282132 476776
rect 219709 476718 282132 476720
rect 219709 476715 219775 476718
rect 282126 476716 282132 476718
rect 282196 476716 282202 476780
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 228541 454066 228607 454069
rect 383929 454066 383995 454069
rect 228541 454064 383995 454066
rect 228541 454008 228546 454064
rect 228602 454008 383934 454064
rect 383990 454008 383995 454064
rect 228541 454006 383995 454008
rect 228541 454003 228607 454006
rect 383929 454003 383995 454006
rect 298001 452434 298067 452437
rect 298001 452432 300196 452434
rect 298001 452376 298006 452432
rect 298062 452376 300196 452432
rect 298001 452374 300196 452376
rect 298001 452371 298067 452374
rect 384021 452298 384087 452301
rect 383886 452296 384087 452298
rect 383886 452240 384026 452296
rect 384082 452240 384087 452296
rect 383886 452238 384087 452240
rect 383886 451724 383946 452238
rect 384021 452235 384087 452238
rect -960 449578 480 449668
rect 2865 449578 2931 449581
rect -960 449576 2931 449578
rect -960 449520 2870 449576
rect 2926 449520 2931 449576
rect -960 449518 2931 449520
rect -960 449428 480 449518
rect 2865 449515 2931 449518
rect 254025 449306 254091 449309
rect 284661 449306 284727 449309
rect 254025 449304 284727 449306
rect 254025 449248 254030 449304
rect 254086 449248 284666 449304
rect 284722 449248 284727 449304
rect 254025 449246 284727 449248
rect 254025 449243 254091 449246
rect 284661 449243 284727 449246
rect 252921 449170 252987 449173
rect 284753 449170 284819 449173
rect 252921 449168 284819 449170
rect 252921 449112 252926 449168
rect 252982 449112 284758 449168
rect 284814 449112 284819 449168
rect 252921 449110 284819 449112
rect 252921 449107 252987 449110
rect 284753 449107 284819 449110
rect 297357 448354 297423 448357
rect 297357 448352 300196 448354
rect 297357 448296 297362 448352
rect 297418 448296 300196 448352
rect 297357 448294 300196 448296
rect 297357 448291 297423 448294
rect 384021 448218 384087 448221
rect 383886 448216 384087 448218
rect 383886 448160 384026 448216
rect 384082 448160 384087 448216
rect 383886 448158 384087 448160
rect 383886 447644 383946 448158
rect 384021 448155 384087 448158
rect 235533 446858 235599 446861
rect 257470 446858 257476 446860
rect 235533 446856 257476 446858
rect 235533 446800 235538 446856
rect 235594 446800 257476 446856
rect 235533 446798 257476 446800
rect 235533 446795 235599 446798
rect 257470 446796 257476 446798
rect 257540 446796 257546 446860
rect 209589 446722 209655 446725
rect 262622 446722 262628 446724
rect 209589 446720 262628 446722
rect 209589 446664 209594 446720
rect 209650 446664 262628 446720
rect 209589 446662 262628 446664
rect 209589 446659 209655 446662
rect 262622 446660 262628 446662
rect 262692 446660 262698 446724
rect 209037 446586 209103 446589
rect 298921 446586 298987 446589
rect 209037 446584 298987 446586
rect 209037 446528 209042 446584
rect 209098 446528 298926 446584
rect 298982 446528 298987 446584
rect 209037 446526 298987 446528
rect 209037 446523 209103 446526
rect 298921 446523 298987 446526
rect 206829 446450 206895 446453
rect 229001 446450 229067 446453
rect 206829 446448 229067 446450
rect 206829 446392 206834 446448
rect 206890 446392 229006 446448
rect 229062 446392 229067 446448
rect 206829 446390 229067 446392
rect 206829 446387 206895 446390
rect 229001 446387 229067 446390
rect 204345 446314 204411 446317
rect 229093 446314 229159 446317
rect 204345 446312 229159 446314
rect 204345 446256 204350 446312
rect 204406 446256 229098 446312
rect 229154 446256 229159 446312
rect 204345 446254 229159 446256
rect 204345 446251 204411 446254
rect 229093 446251 229159 446254
rect 233601 446314 233667 446317
rect 264421 446314 264487 446317
rect 233601 446312 264487 446314
rect 233601 446256 233606 446312
rect 233662 446256 264426 446312
rect 264482 446256 264487 446312
rect 233601 446254 264487 446256
rect 233601 446251 233667 446254
rect 264421 446251 264487 446254
rect 204621 446178 204687 446181
rect 229737 446178 229803 446181
rect 204621 446176 229803 446178
rect 204621 446120 204626 446176
rect 204682 446120 229742 446176
rect 229798 446120 229803 446176
rect 204621 446118 229803 446120
rect 204621 446115 204687 446118
rect 229737 446115 229803 446118
rect 237741 446178 237807 446181
rect 254526 446178 254532 446180
rect 237741 446176 254532 446178
rect 237741 446120 237746 446176
rect 237802 446120 254532 446176
rect 237741 446118 254532 446120
rect 237741 446115 237807 446118
rect 254526 446116 254532 446118
rect 254596 446116 254602 446180
rect 260833 446178 260899 446181
rect 298502 446178 298508 446180
rect 260833 446176 298508 446178
rect 260833 446120 260838 446176
rect 260894 446120 298508 446176
rect 260833 446118 298508 446120
rect 260833 446115 260899 446118
rect 298502 446116 298508 446118
rect 298572 446116 298578 446180
rect 201953 446042 202019 446045
rect 234705 446042 234771 446045
rect 201953 446040 234771 446042
rect 201953 445984 201958 446040
rect 202014 445984 234710 446040
rect 234766 445984 234771 446040
rect 201953 445982 234771 445984
rect 201953 445979 202019 445982
rect 234705 445979 234771 445982
rect 251725 446042 251791 446045
rect 296069 446042 296135 446045
rect 251725 446040 296135 446042
rect 251725 445984 251730 446040
rect 251786 445984 296074 446040
rect 296130 445984 296135 446040
rect 251725 445982 296135 445984
rect 251725 445979 251791 445982
rect 296069 445979 296135 445982
rect 251817 445906 251883 445909
rect 265801 445906 265867 445909
rect 251817 445904 265867 445906
rect 251817 445848 251822 445904
rect 251878 445848 265806 445904
rect 265862 445848 265867 445904
rect 251817 445846 265867 445848
rect 251817 445843 251883 445846
rect 265801 445843 265867 445846
rect 250437 445770 250503 445773
rect 257286 445770 257292 445772
rect 250437 445768 257292 445770
rect 250437 445712 250442 445768
rect 250498 445712 257292 445768
rect 250437 445710 257292 445712
rect 250437 445707 250503 445710
rect 257286 445708 257292 445710
rect 257356 445708 257362 445772
rect 245469 445634 245535 445637
rect 254894 445634 254900 445636
rect 245469 445632 254900 445634
rect 245469 445576 245474 445632
rect 245530 445576 254900 445632
rect 245469 445574 254900 445576
rect 245469 445571 245535 445574
rect 254894 445572 254900 445574
rect 254964 445572 254970 445636
rect 258441 445634 258507 445637
rect 260598 445634 260604 445636
rect 258441 445632 260604 445634
rect 258441 445576 258446 445632
rect 258502 445576 260604 445632
rect 258441 445574 260604 445576
rect 258441 445571 258507 445574
rect 260598 445572 260604 445574
rect 260668 445572 260674 445636
rect 235257 445090 235323 445093
rect 254710 445090 254716 445092
rect 235257 445088 254716 445090
rect 235257 445032 235262 445088
rect 235318 445032 254716 445088
rect 235257 445030 254716 445032
rect 235257 445027 235323 445030
rect 254710 445028 254716 445030
rect 254780 445028 254786 445092
rect 207105 444954 207171 444957
rect 272517 444954 272583 444957
rect 207105 444952 272583 444954
rect 207105 444896 207110 444952
rect 207166 444896 272522 444952
rect 272578 444896 272583 444952
rect 207105 444894 272583 444896
rect 207105 444891 207171 444894
rect 272517 444891 272583 444894
rect 205449 444818 205515 444821
rect 264237 444818 264303 444821
rect 205449 444816 264303 444818
rect 205449 444760 205454 444816
rect 205510 444760 264242 444816
rect 264298 444760 264303 444816
rect 205449 444758 264303 444760
rect 205449 444755 205515 444758
rect 264237 444755 264303 444758
rect 205725 444682 205791 444685
rect 265709 444682 265775 444685
rect 205725 444680 265775 444682
rect 205725 444624 205730 444680
rect 205786 444624 265714 444680
rect 265770 444624 265775 444680
rect 583520 444668 584960 444908
rect 205725 444622 265775 444624
rect 205725 444619 205791 444622
rect 265709 444619 265775 444622
rect 206277 444546 206343 444549
rect 266997 444546 267063 444549
rect 206277 444544 267063 444546
rect 206277 444488 206282 444544
rect 206338 444488 267002 444544
rect 267058 444488 267063 444544
rect 206277 444486 267063 444488
rect 206277 444483 206343 444486
rect 266997 444483 267063 444486
rect 251541 444410 251607 444413
rect 260046 444410 260052 444412
rect 251541 444408 260052 444410
rect 251541 444352 251546 444408
rect 251602 444352 260052 444408
rect 251541 444350 260052 444352
rect 251541 444347 251607 444350
rect 260046 444348 260052 444350
rect 260116 444348 260122 444412
rect 213085 444138 213151 444141
rect 247493 444138 247559 444141
rect 253790 444138 253796 444140
rect 213085 444136 218070 444138
rect 213085 444080 213090 444136
rect 213146 444080 218070 444136
rect 213085 444078 218070 444080
rect 213085 444075 213151 444078
rect 217409 444002 217475 444005
rect 208350 444000 217475 444002
rect 208350 443944 217414 444000
rect 217470 443944 217475 444000
rect 208350 443942 217475 443944
rect 218010 444002 218070 444078
rect 247493 444136 253796 444138
rect 247493 444080 247498 444136
rect 247554 444080 253796 444136
rect 247493 444078 253796 444080
rect 247493 444075 247559 444078
rect 253790 444076 253796 444078
rect 253860 444076 253866 444140
rect 220445 444002 220511 444005
rect 218010 444000 220511 444002
rect 218010 443944 220450 444000
rect 220506 443944 220511 444000
rect 218010 443942 220511 443944
rect 207565 443866 207631 443869
rect 208350 443866 208410 443942
rect 217409 443939 217475 443942
rect 220445 443939 220511 443942
rect 207565 443864 208410 443866
rect 207565 443808 207570 443864
rect 207626 443808 208410 443864
rect 207565 443806 208410 443808
rect 211061 443866 211127 443869
rect 212942 443866 212948 443868
rect 211061 443864 212948 443866
rect 211061 443808 211066 443864
rect 211122 443808 212948 443864
rect 211061 443806 212948 443808
rect 207565 443803 207631 443806
rect 211061 443803 211127 443806
rect 212942 443804 212948 443806
rect 213012 443804 213018 443868
rect 219341 443866 219407 443869
rect 232313 443868 232379 443869
rect 233233 443868 233299 443869
rect 234889 443868 234955 443869
rect 232262 443866 232268 443868
rect 213134 443864 219407 443866
rect 213134 443808 219346 443864
rect 219402 443808 219407 443864
rect 213134 443806 219407 443808
rect 232222 443806 232268 443866
rect 232332 443864 232379 443868
rect 233182 443866 233188 443868
rect 232374 443808 232379 443864
rect 203425 443730 203491 443733
rect 213134 443730 213194 443806
rect 219341 443803 219407 443806
rect 232262 443804 232268 443806
rect 232332 443804 232379 443808
rect 233142 443806 233188 443866
rect 233252 443864 233299 443868
rect 234838 443866 234844 443868
rect 233294 443808 233299 443864
rect 233182 443804 233188 443806
rect 233252 443804 233299 443808
rect 234798 443806 234844 443866
rect 234908 443864 234955 443868
rect 234950 443808 234955 443864
rect 234838 443804 234844 443806
rect 234908 443804 234955 443808
rect 232313 443803 232379 443804
rect 233233 443803 233299 443804
rect 234889 443803 234955 443804
rect 203425 443728 213194 443730
rect 203425 443672 203430 443728
rect 203486 443672 213194 443728
rect 203425 443670 213194 443672
rect 217409 443730 217475 443733
rect 298737 443730 298803 443733
rect 217409 443728 298803 443730
rect 217409 443672 217414 443728
rect 217470 443672 298742 443728
rect 298798 443672 298803 443728
rect 217409 443670 298803 443672
rect 203425 443667 203491 443670
rect 217409 443667 217475 443670
rect 298737 443667 298803 443670
rect 205081 443594 205147 443597
rect 256601 443596 256667 443597
rect 205081 443592 213194 443594
rect 205081 443536 205086 443592
rect 205142 443536 213194 443592
rect 205081 443534 213194 443536
rect 205081 443531 205147 443534
rect 205357 443458 205423 443461
rect 206185 443458 206251 443461
rect 210366 443458 210372 443460
rect 205357 443456 205650 443458
rect 205357 443400 205362 443456
rect 205418 443400 205650 443456
rect 205357 443398 205650 443400
rect 205357 443395 205423 443398
rect 205590 443186 205650 443398
rect 206185 443456 210372 443458
rect 206185 443400 206190 443456
rect 206246 443400 210372 443456
rect 206185 443398 210372 443400
rect 206185 443395 206251 443398
rect 210366 443396 210372 443398
rect 210436 443396 210442 443460
rect 210601 443458 210667 443461
rect 213134 443458 213194 443534
rect 214230 443532 214236 443596
rect 214300 443594 214306 443596
rect 255814 443594 255820 443596
rect 214300 443534 255820 443594
rect 214300 443532 214306 443534
rect 255814 443532 255820 443534
rect 255884 443532 255890 443596
rect 256550 443594 256556 443596
rect 256510 443534 256556 443594
rect 256620 443592 256667 443596
rect 265617 443594 265683 443597
rect 256662 443536 256667 443592
rect 256550 443532 256556 443534
rect 256620 443532 256667 443536
rect 256601 443531 256667 443532
rect 258766 443592 265683 443594
rect 258766 443536 265622 443592
rect 265678 443536 265683 443592
rect 258766 443534 265683 443536
rect 258766 443458 258826 443534
rect 265617 443531 265683 443534
rect 298001 443594 298067 443597
rect 298001 443592 300196 443594
rect 298001 443536 298006 443592
rect 298062 443536 300196 443592
rect 298001 443534 300196 443536
rect 298001 443531 298067 443534
rect 210601 443456 213010 443458
rect 210601 443400 210606 443456
rect 210662 443400 213010 443456
rect 210601 443398 213010 443400
rect 213134 443398 258826 443458
rect 258901 443458 258967 443461
rect 259361 443460 259427 443461
rect 262121 443460 262187 443461
rect 259126 443458 259132 443460
rect 258901 443456 259132 443458
rect 258901 443400 258906 443456
rect 258962 443400 259132 443456
rect 258901 443398 259132 443400
rect 210601 443395 210667 443398
rect 212950 443322 213010 443398
rect 258901 443395 258967 443398
rect 259126 443396 259132 443398
rect 259196 443396 259202 443460
rect 259310 443458 259316 443460
rect 259270 443398 259316 443458
rect 259380 443456 259427 443460
rect 262070 443458 262076 443460
rect 259422 443400 259427 443456
rect 259310 443396 259316 443398
rect 259380 443396 259427 443400
rect 262030 443398 262076 443458
rect 262140 443456 262187 443460
rect 262182 443400 262187 443456
rect 262070 443396 262076 443398
rect 262140 443396 262187 443400
rect 259361 443395 259427 443396
rect 262121 443395 262187 443396
rect 214230 443322 214236 443324
rect 212950 443262 214236 443322
rect 214230 443260 214236 443262
rect 214300 443260 214306 443324
rect 214414 443260 214420 443324
rect 214484 443322 214490 443324
rect 296161 443322 296227 443325
rect 214484 443320 296227 443322
rect 214484 443264 296166 443320
rect 296222 443264 296227 443320
rect 214484 443262 296227 443264
rect 214484 443260 214490 443262
rect 296161 443259 296227 443262
rect 295977 443186 296043 443189
rect 205590 443184 296043 443186
rect 205590 443128 295982 443184
rect 296038 443128 296043 443184
rect 205590 443126 296043 443128
rect 295977 443123 296043 443126
rect 210366 442988 210372 443052
rect 210436 443050 210442 443052
rect 214414 443050 214420 443052
rect 210436 442990 214420 443050
rect 210436 442988 210442 442990
rect 214414 442988 214420 442990
rect 214484 442988 214490 443052
rect 385493 442914 385559 442917
rect 383916 442912 385559 442914
rect 383916 442856 385498 442912
rect 385554 442856 385559 442912
rect 383916 442854 385559 442856
rect 385493 442851 385559 442854
rect 202689 442642 202755 442645
rect 232262 442642 232268 442644
rect 202689 442640 232268 442642
rect 202689 442584 202694 442640
rect 202750 442584 232268 442640
rect 202689 442582 232268 442584
rect 202689 442579 202755 442582
rect 232262 442580 232268 442582
rect 232332 442580 232338 442644
rect 202505 442506 202571 442509
rect 233182 442506 233188 442508
rect 202505 442504 233188 442506
rect 202505 442448 202510 442504
rect 202566 442448 233188 442504
rect 202505 442446 233188 442448
rect 202505 442443 202571 442446
rect 233182 442444 233188 442446
rect 233252 442444 233258 442508
rect 202137 442370 202203 442373
rect 234838 442370 234844 442372
rect 202137 442368 234844 442370
rect 202137 442312 202142 442368
rect 202198 442312 234844 442368
rect 202137 442310 234844 442312
rect 202137 442307 202203 442310
rect 234838 442308 234844 442310
rect 234908 442308 234914 442372
rect 212942 442172 212948 442236
rect 213012 442234 213018 442236
rect 296621 442234 296687 442237
rect 213012 442232 296687 442234
rect 213012 442176 296626 442232
rect 296682 442176 296687 442232
rect 213012 442174 296687 442176
rect 213012 442172 213018 442174
rect 296621 442171 296687 442174
rect 298001 439514 298067 439517
rect 298001 439512 300196 439514
rect 298001 439456 298006 439512
rect 298062 439456 300196 439512
rect 298001 439454 300196 439456
rect 298001 439451 298067 439454
rect 383886 438701 383946 438804
rect 383886 438696 383995 438701
rect 383886 438640 383934 438696
rect 383990 438640 383995 438696
rect 383886 438638 383995 438640
rect 383929 438635 383995 438638
rect -960 436508 480 436748
rect 298001 434754 298067 434757
rect 298001 434752 300196 434754
rect 298001 434696 298006 434752
rect 298062 434696 300196 434752
rect 298001 434694 300196 434696
rect 298001 434691 298067 434694
rect 385401 434074 385467 434077
rect 383916 434072 385467 434074
rect 383916 434016 385406 434072
rect 385462 434016 385467 434072
rect 383916 434014 385467 434016
rect 385401 434011 385467 434014
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 298001 430674 298067 430677
rect 298001 430672 300196 430674
rect 298001 430616 298006 430672
rect 298062 430616 300196 430672
rect 298001 430614 300196 430616
rect 298001 430611 298067 430614
rect 385309 429994 385375 429997
rect 383916 429992 385375 429994
rect 383916 429936 385314 429992
rect 385370 429936 385375 429992
rect 383916 429934 385375 429936
rect 385309 429931 385375 429934
rect 298001 425914 298067 425917
rect 298001 425912 300196 425914
rect 298001 425856 298006 425912
rect 298062 425856 300196 425912
rect 298001 425854 300196 425856
rect 298001 425851 298067 425854
rect 385217 425234 385283 425237
rect 383916 425232 385283 425234
rect 383916 425176 385222 425232
rect 385278 425176 385283 425232
rect 383916 425174 385283 425176
rect 385217 425171 385283 425174
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 297909 421834 297975 421837
rect 297909 421832 300196 421834
rect 297909 421776 297914 421832
rect 297970 421776 300196 421832
rect 297909 421774 300196 421776
rect 297909 421771 297975 421774
rect 383929 421698 383995 421701
rect 383886 421696 383995 421698
rect 383886 421640 383934 421696
rect 383990 421640 383995 421696
rect 383886 421635 383995 421640
rect 383886 421124 383946 421635
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 297633 417074 297699 417077
rect 297633 417072 300196 417074
rect 297633 417016 297638 417072
rect 297694 417016 300196 417072
rect 297633 417014 300196 417016
rect 297633 417011 297699 417014
rect 385125 416394 385191 416397
rect 383916 416392 385191 416394
rect 383916 416336 385130 416392
rect 385186 416336 385191 416392
rect 383916 416334 385191 416336
rect 385125 416331 385191 416334
rect 297541 412994 297607 412997
rect 297541 412992 300196 412994
rect 297541 412936 297546 412992
rect 297602 412936 300196 412992
rect 297541 412934 300196 412936
rect 297541 412931 297607 412934
rect 385033 412314 385099 412317
rect 383916 412312 385099 412314
rect 383916 412256 385038 412312
rect 385094 412256 385099 412312
rect 383916 412254 385099 412256
rect 385033 412251 385099 412254
rect -960 410546 480 410636
rect 3509 410546 3575 410549
rect -960 410544 3575 410546
rect -960 410488 3514 410544
rect 3570 410488 3575 410544
rect -960 410486 3575 410488
rect -960 410396 480 410486
rect 3509 410483 3575 410486
rect 298001 408234 298067 408237
rect 298001 408232 300196 408234
rect 298001 408176 298006 408232
rect 298062 408176 300196 408232
rect 298001 408174 300196 408176
rect 298001 408171 298067 408174
rect 385033 407554 385099 407557
rect 383916 407552 385099 407554
rect 383916 407496 385038 407552
rect 385094 407496 385099 407552
rect 383916 407494 385099 407496
rect 385033 407491 385099 407494
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect 296989 404154 297055 404157
rect 296989 404152 300196 404154
rect 296989 404096 296994 404152
rect 297050 404096 300196 404152
rect 296989 404094 300196 404096
rect 296989 404091 297055 404094
rect 383334 402932 383394 403444
rect 383326 402868 383332 402932
rect 383396 402868 383402 402932
rect 259126 401508 259132 401572
rect 259196 401570 259202 401572
rect 383326 401570 383332 401572
rect 259196 401510 383332 401570
rect 259196 401508 259202 401510
rect 383326 401508 383332 401510
rect 383396 401508 383402 401572
rect 256550 400148 256556 400212
rect 256620 400210 256626 400212
rect 260005 400210 260071 400213
rect 256620 400208 260071 400210
rect 256620 400152 260010 400208
rect 260066 400152 260071 400208
rect 256620 400150 260071 400152
rect 256620 400148 256626 400150
rect 260005 400147 260071 400150
rect 253054 399468 253060 399532
rect 253124 399530 253130 399532
rect 253657 399530 253723 399533
rect 253124 399528 253723 399530
rect 253124 399472 253662 399528
rect 253718 399472 253723 399528
rect 253124 399470 253723 399472
rect 253124 399468 253130 399470
rect 253657 399467 253723 399470
rect 253790 399468 253796 399532
rect 253860 399530 253866 399532
rect 580257 399530 580323 399533
rect 253860 399528 580323 399530
rect 253860 399472 580262 399528
rect 580318 399472 580323 399528
rect 253860 399470 580323 399472
rect 253860 399468 253866 399470
rect 580257 399467 580323 399470
rect 253105 399394 253171 399397
rect 253238 399394 253244 399396
rect 253105 399392 253244 399394
rect 253105 399336 253110 399392
rect 253166 399336 253244 399392
rect 253105 399334 253244 399336
rect 253105 399331 253171 399334
rect 253238 399332 253244 399334
rect 253308 399332 253314 399396
rect 255221 399260 255287 399261
rect 255221 399256 255268 399260
rect 255332 399258 255338 399260
rect 255221 399200 255226 399256
rect 255221 399196 255268 399200
rect 255332 399198 255378 399258
rect 255332 399196 255338 399198
rect 255221 399195 255287 399196
rect 245377 399122 245443 399125
rect 245377 399120 253950 399122
rect 245377 399064 245382 399120
rect 245438 399064 253950 399120
rect 245377 399062 253950 399064
rect 245377 399059 245443 399062
rect 216765 398986 216831 398989
rect 242801 398986 242867 398989
rect 216765 398984 216874 398986
rect 216765 398928 216770 398984
rect 216826 398928 216874 398984
rect 216765 398923 216874 398928
rect 208209 398850 208275 398853
rect 212165 398850 212231 398853
rect 208209 398848 212231 398850
rect 208209 398792 208214 398848
rect 208270 398792 212170 398848
rect 212226 398792 212231 398848
rect 208209 398790 212231 398792
rect 216814 398850 216874 398923
rect 242758 398984 242867 398986
rect 242758 398928 242806 398984
rect 242862 398928 242867 398984
rect 242758 398923 242867 398928
rect 217174 398850 217180 398852
rect 216814 398790 217180 398850
rect 208209 398787 208275 398790
rect 212165 398787 212231 398790
rect 217174 398788 217180 398790
rect 217244 398788 217250 398852
rect 207749 398714 207815 398717
rect 212625 398714 212691 398717
rect 207749 398712 212691 398714
rect 207749 398656 207754 398712
rect 207810 398656 212630 398712
rect 212686 398656 212691 398712
rect 207749 398654 212691 398656
rect 207749 398651 207815 398654
rect 212625 398651 212691 398654
rect 242617 398714 242683 398717
rect 242758 398714 242818 398923
rect 242617 398712 242818 398714
rect 242617 398656 242622 398712
rect 242678 398656 242818 398712
rect 242617 398654 242818 398656
rect 253197 398716 253263 398717
rect 253197 398712 253244 398716
rect 253308 398714 253314 398716
rect 253890 398714 253950 399062
rect 254526 399060 254532 399124
rect 254596 399122 254602 399124
rect 257245 399122 257311 399125
rect 254596 399120 257311 399122
rect 254596 399064 257250 399120
rect 257306 399064 257311 399120
rect 254596 399062 257311 399064
rect 254596 399060 254602 399062
rect 257245 399059 257311 399062
rect 257470 399060 257476 399124
rect 257540 399122 257546 399124
rect 312261 399122 312327 399125
rect 324497 399122 324563 399125
rect 257540 399120 312327 399122
rect 257540 399064 312266 399120
rect 312322 399064 312327 399120
rect 257540 399062 312327 399064
rect 257540 399060 257546 399062
rect 312261 399059 312327 399062
rect 321510 399120 324563 399122
rect 321510 399064 324502 399120
rect 324558 399064 324563 399120
rect 321510 399062 324563 399064
rect 254894 398924 254900 398988
rect 254964 398986 254970 398988
rect 321510 398986 321570 399062
rect 324497 399059 324563 399062
rect 254964 398926 321570 398986
rect 321694 398926 331230 398986
rect 254964 398924 254970 398926
rect 321694 398850 321754 398926
rect 263366 398790 321754 398850
rect 331170 398850 331230 398926
rect 379237 398850 379303 398853
rect 331170 398848 379303 398850
rect 331170 398792 379242 398848
rect 379298 398792 379303 398848
rect 331170 398790 379303 398792
rect 257245 398714 257311 398717
rect 263366 398714 263426 398790
rect 379237 398787 379303 398790
rect 253197 398656 253202 398712
rect 242617 398651 242683 398654
rect 253197 398652 253244 398656
rect 253308 398654 253354 398714
rect 253890 398654 256434 398714
rect 253308 398652 253314 398654
rect 253197 398651 253263 398652
rect 206277 398578 206343 398581
rect 212809 398578 212875 398581
rect 206277 398576 212875 398578
rect 206277 398520 206282 398576
rect 206338 398520 212814 398576
rect 212870 398520 212875 398576
rect 206277 398518 212875 398520
rect 206277 398515 206343 398518
rect 212809 398515 212875 398518
rect 248781 398578 248847 398581
rect 256233 398578 256299 398581
rect 248781 398576 256299 398578
rect 248781 398520 248786 398576
rect 248842 398520 256238 398576
rect 256294 398520 256299 398576
rect 248781 398518 256299 398520
rect 256374 398578 256434 398654
rect 257245 398712 263426 398714
rect 257245 398656 257250 398712
rect 257306 398656 263426 398712
rect 257245 398654 263426 398656
rect 263501 398714 263567 398717
rect 362493 398714 362559 398717
rect 263501 398712 362559 398714
rect 263501 398656 263506 398712
rect 263562 398656 362498 398712
rect 362554 398656 362559 398712
rect 263501 398654 362559 398656
rect 257245 398651 257311 398654
rect 263501 398651 263567 398654
rect 362493 398651 362559 398654
rect 258809 398578 258875 398581
rect 256374 398576 258875 398578
rect 256374 398520 258814 398576
rect 258870 398520 258875 398576
rect 256374 398518 258875 398520
rect 248781 398515 248847 398518
rect 256233 398515 256299 398518
rect 258809 398515 258875 398518
rect 260046 398516 260052 398580
rect 260116 398578 260122 398580
rect 357985 398578 358051 398581
rect 260116 398576 358051 398578
rect 260116 398520 357990 398576
rect 358046 398520 358051 398576
rect 260116 398518 358051 398520
rect 260116 398516 260122 398518
rect 357985 398515 358051 398518
rect 211521 398442 211587 398445
rect 219341 398442 219407 398445
rect 200070 398440 211587 398442
rect 200070 398384 211526 398440
rect 211582 398384 211587 398440
rect 200070 398382 211587 398384
rect 42057 398034 42123 398037
rect 200070 398034 200130 398382
rect 211521 398379 211587 398382
rect 219206 398440 219407 398442
rect 219206 398384 219346 398440
rect 219402 398384 219407 398440
rect 219206 398382 219407 398384
rect 210233 398170 210299 398173
rect 213913 398170 213979 398173
rect 210233 398168 213979 398170
rect 210233 398112 210238 398168
rect 210294 398112 213918 398168
rect 213974 398112 213979 398168
rect 210233 398110 213979 398112
rect 210233 398107 210299 398110
rect 213913 398107 213979 398110
rect 213361 398034 213427 398037
rect 215293 398034 215359 398037
rect 42057 398032 200130 398034
rect 42057 397976 42062 398032
rect 42118 397976 200130 398032
rect 42057 397974 200130 397976
rect 210558 398032 213427 398034
rect 210558 397976 213366 398032
rect 213422 397976 213427 398032
rect 210558 397974 213427 397976
rect 42057 397971 42123 397974
rect 209814 397700 209820 397764
rect 209884 397762 209890 397764
rect 210325 397762 210391 397765
rect 209884 397760 210391 397762
rect 209884 397704 210330 397760
rect 210386 397704 210391 397760
rect 209884 397702 210391 397704
rect 209884 397700 209890 397702
rect 210325 397699 210391 397702
rect 204989 397626 205055 397629
rect 210233 397626 210299 397629
rect 204989 397624 210299 397626
rect -960 397490 480 397580
rect 204989 397568 204994 397624
rect 205050 397568 210238 397624
rect 210294 397568 210299 397624
rect 204989 397566 210299 397568
rect 204989 397563 205055 397566
rect 210233 397563 210299 397566
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 206461 397490 206527 397493
rect 210558 397490 210618 397974
rect 213361 397971 213427 397974
rect 213502 398032 215359 398034
rect 213502 397976 215298 398032
rect 215354 397976 215359 398032
rect 213502 397974 215359 397976
rect 210693 397898 210759 397901
rect 211429 397898 211495 397901
rect 210693 397896 211495 397898
rect 210693 397840 210698 397896
rect 210754 397840 211434 397896
rect 211490 397840 211495 397896
rect 210693 397838 211495 397840
rect 210693 397835 210759 397838
rect 211429 397835 211495 397838
rect 212625 397898 212691 397901
rect 213502 397898 213562 397974
rect 215293 397971 215359 397974
rect 212625 397896 213562 397898
rect 212625 397840 212630 397896
rect 212686 397840 213562 397896
rect 212625 397838 213562 397840
rect 214005 397898 214071 397901
rect 214414 397898 214420 397900
rect 214005 397896 214420 397898
rect 214005 397840 214010 397896
rect 214066 397840 214420 397896
rect 214005 397838 214420 397840
rect 212625 397835 212691 397838
rect 214005 397835 214071 397838
rect 214414 397836 214420 397838
rect 214484 397836 214490 397900
rect 217133 397898 217199 397901
rect 214974 397896 217199 397898
rect 214974 397840 217138 397896
rect 217194 397840 217199 397896
rect 214974 397838 217199 397840
rect 211102 397700 211108 397764
rect 211172 397762 211178 397764
rect 211613 397762 211679 397765
rect 211172 397760 211679 397762
rect 211172 397704 211618 397760
rect 211674 397704 211679 397760
rect 211172 397702 211679 397704
rect 211172 397700 211178 397702
rect 211613 397699 211679 397702
rect 212257 397762 212323 397765
rect 214741 397762 214807 397765
rect 212257 397760 214807 397762
rect 212257 397704 212262 397760
rect 212318 397704 214746 397760
rect 214802 397704 214807 397760
rect 212257 397702 214807 397704
rect 212257 397699 212323 397702
rect 214741 397699 214807 397702
rect 211245 397626 211311 397629
rect 211470 397626 211476 397628
rect 211245 397624 211476 397626
rect 211245 397568 211250 397624
rect 211306 397568 211476 397624
rect 211245 397566 211476 397568
rect 211245 397563 211311 397566
rect 211470 397564 211476 397566
rect 211540 397564 211546 397628
rect 214046 397564 214052 397628
rect 214116 397626 214122 397628
rect 214281 397626 214347 397629
rect 214116 397624 214347 397626
rect 214116 397568 214286 397624
rect 214342 397568 214347 397624
rect 214116 397566 214347 397568
rect 214116 397564 214122 397566
rect 214281 397563 214347 397566
rect 214741 397626 214807 397629
rect 214974 397626 215034 397838
rect 217133 397835 217199 397838
rect 218881 397898 218947 397901
rect 219206 397898 219266 398382
rect 219341 398379 219407 398382
rect 247309 398442 247375 398445
rect 253657 398442 253723 398445
rect 247309 398440 253723 398442
rect 247309 398384 247314 398440
rect 247370 398384 253662 398440
rect 253718 398384 253723 398440
rect 247309 398382 253723 398384
rect 247309 398379 247375 398382
rect 253657 398379 253723 398382
rect 257286 398380 257292 398444
rect 257356 398442 257362 398444
rect 263409 398442 263475 398445
rect 257356 398440 263475 398442
rect 257356 398384 263414 398440
rect 263470 398384 263475 398440
rect 257356 398382 263475 398384
rect 257356 398380 257362 398382
rect 263409 398379 263475 398382
rect 263542 398380 263548 398444
rect 263612 398442 263618 398444
rect 332869 398442 332935 398445
rect 263612 398440 332935 398442
rect 263612 398384 332874 398440
rect 332930 398384 332935 398440
rect 263612 398382 332935 398384
rect 263612 398380 263618 398382
rect 332869 398379 332935 398382
rect 219341 398306 219407 398309
rect 219801 398306 219867 398309
rect 219341 398304 219867 398306
rect 219341 398248 219346 398304
rect 219402 398248 219806 398304
rect 219862 398248 219867 398304
rect 219341 398246 219867 398248
rect 219341 398243 219407 398246
rect 219801 398243 219867 398246
rect 251265 398306 251331 398309
rect 253105 398306 253171 398309
rect 251265 398304 253171 398306
rect 251265 398248 251270 398304
rect 251326 398248 253110 398304
rect 253166 398248 253171 398304
rect 251265 398246 253171 398248
rect 251265 398243 251331 398246
rect 253105 398243 253171 398246
rect 255589 398306 255655 398309
rect 256785 398306 256851 398309
rect 255589 398304 256851 398306
rect 255589 398248 255594 398304
rect 255650 398248 256790 398304
rect 256846 398248 256851 398304
rect 255589 398246 256851 398248
rect 255589 398243 255655 398246
rect 256785 398243 256851 398246
rect 259310 398244 259316 398308
rect 259380 398306 259386 398308
rect 316125 398306 316191 398309
rect 259380 398304 316191 398306
rect 259380 398248 316130 398304
rect 316186 398248 316191 398304
rect 259380 398246 316191 398248
rect 259380 398244 259386 398246
rect 316125 398243 316191 398246
rect 248505 398170 248571 398173
rect 489913 398170 489979 398173
rect 248505 398168 489979 398170
rect 248505 398112 248510 398168
rect 248566 398112 489918 398168
rect 489974 398112 489979 398168
rect 248505 398110 489979 398112
rect 248505 398107 248571 398110
rect 489913 398107 489979 398110
rect 226190 397972 226196 398036
rect 226260 398034 226266 398036
rect 233601 398034 233667 398037
rect 226260 398032 233667 398034
rect 226260 397976 233606 398032
rect 233662 397976 233667 398032
rect 226260 397974 233667 397976
rect 226260 397972 226266 397974
rect 233601 397971 233667 397974
rect 249885 398034 249951 398037
rect 507853 398034 507919 398037
rect 249885 398032 507919 398034
rect 249885 397976 249890 398032
rect 249946 397976 507858 398032
rect 507914 397976 507919 398032
rect 249885 397974 507919 397976
rect 249885 397971 249951 397974
rect 507853 397971 507919 397974
rect 218881 397896 219266 397898
rect 218881 397840 218886 397896
rect 218942 397840 219266 397896
rect 218881 397838 219266 397840
rect 223757 397898 223823 397901
rect 224166 397898 224172 397900
rect 223757 397896 224172 397898
rect 223757 397840 223762 397896
rect 223818 397840 224172 397896
rect 223757 397838 224172 397840
rect 218881 397835 218947 397838
rect 223757 397835 223823 397838
rect 224166 397836 224172 397838
rect 224236 397836 224242 397900
rect 230197 397898 230263 397901
rect 230422 397898 230428 397900
rect 230197 397896 230428 397898
rect 230197 397840 230202 397896
rect 230258 397840 230428 397896
rect 230197 397838 230428 397840
rect 230197 397835 230263 397838
rect 230422 397836 230428 397838
rect 230492 397836 230498 397900
rect 239438 397836 239444 397900
rect 239508 397898 239514 397900
rect 240041 397898 240107 397901
rect 239508 397896 240107 397898
rect 239508 397840 240046 397896
rect 240102 397840 240107 397896
rect 239508 397838 240107 397840
rect 239508 397836 239514 397838
rect 240041 397835 240107 397838
rect 243486 397836 243492 397900
rect 243556 397898 243562 397900
rect 243905 397898 243971 397901
rect 243556 397896 243971 397898
rect 243556 397840 243910 397896
rect 243966 397840 243971 397896
rect 243556 397838 243971 397840
rect 243556 397836 243562 397838
rect 243905 397835 243971 397838
rect 250897 397898 250963 397901
rect 251030 397898 251036 397900
rect 250897 397896 251036 397898
rect 250897 397840 250902 397896
rect 250958 397840 251036 397896
rect 250897 397838 251036 397840
rect 250897 397835 250963 397838
rect 251030 397836 251036 397838
rect 251100 397836 251106 397900
rect 251766 397836 251772 397900
rect 251836 397898 251842 397900
rect 252461 397898 252527 397901
rect 251836 397896 252527 397898
rect 251836 397840 252466 397896
rect 252522 397840 252527 397896
rect 251836 397838 252527 397840
rect 251836 397836 251842 397838
rect 252461 397835 252527 397838
rect 253657 397898 253723 397901
rect 253657 397896 253950 397898
rect 253657 397840 253662 397896
rect 253718 397840 253950 397896
rect 253657 397838 253950 397840
rect 253657 397835 253723 397838
rect 215569 397762 215635 397765
rect 215886 397762 215892 397764
rect 215569 397760 215892 397762
rect 215569 397704 215574 397760
rect 215630 397704 215892 397760
rect 215569 397702 215892 397704
rect 215569 397699 215635 397702
rect 215886 397700 215892 397702
rect 215956 397700 215962 397764
rect 216673 397762 216739 397765
rect 216990 397762 216996 397764
rect 216673 397760 216996 397762
rect 216673 397704 216678 397760
rect 216734 397704 216996 397760
rect 216673 397702 216996 397704
rect 216673 397699 216739 397702
rect 216990 397700 216996 397702
rect 217060 397700 217066 397764
rect 218053 397762 218119 397765
rect 219014 397762 219020 397764
rect 218053 397760 219020 397762
rect 218053 397704 218058 397760
rect 218114 397704 219020 397760
rect 218053 397702 219020 397704
rect 218053 397699 218119 397702
rect 219014 397700 219020 397702
rect 219084 397700 219090 397764
rect 219617 397762 219683 397765
rect 219750 397762 219756 397764
rect 219617 397760 219756 397762
rect 219617 397704 219622 397760
rect 219678 397704 219756 397760
rect 219617 397702 219756 397704
rect 219617 397699 219683 397702
rect 219750 397700 219756 397702
rect 219820 397700 219826 397764
rect 220813 397762 220879 397765
rect 221222 397762 221228 397764
rect 220813 397760 221228 397762
rect 220813 397704 220818 397760
rect 220874 397704 221228 397760
rect 220813 397702 221228 397704
rect 220813 397699 220879 397702
rect 221222 397700 221228 397702
rect 221292 397700 221298 397764
rect 223614 397700 223620 397764
rect 223684 397762 223690 397764
rect 223941 397762 224007 397765
rect 223684 397760 224007 397762
rect 223684 397704 223946 397760
rect 224002 397704 224007 397760
rect 223684 397702 224007 397704
rect 223684 397700 223690 397702
rect 223941 397699 224007 397702
rect 228582 397700 228588 397764
rect 228652 397762 228658 397764
rect 228817 397762 228883 397765
rect 228652 397760 228883 397762
rect 228652 397704 228822 397760
rect 228878 397704 228883 397760
rect 228652 397702 228883 397704
rect 228652 397700 228658 397702
rect 228817 397699 228883 397702
rect 229870 397700 229876 397764
rect 229940 397762 229946 397764
rect 230289 397762 230355 397765
rect 229940 397760 230355 397762
rect 229940 397704 230294 397760
rect 230350 397704 230355 397760
rect 229940 397702 230355 397704
rect 229940 397700 229946 397702
rect 230289 397699 230355 397702
rect 232630 397700 232636 397764
rect 232700 397762 232706 397764
rect 232957 397762 233023 397765
rect 232700 397760 233023 397762
rect 232700 397704 232962 397760
rect 233018 397704 233023 397760
rect 232700 397702 233023 397704
rect 232700 397700 232706 397702
rect 232957 397699 233023 397702
rect 233918 397700 233924 397764
rect 233988 397762 233994 397764
rect 234429 397762 234495 397765
rect 233988 397760 234495 397762
rect 233988 397704 234434 397760
rect 234490 397704 234495 397760
rect 233988 397702 234495 397704
rect 233988 397700 233994 397702
rect 234429 397699 234495 397702
rect 236862 397700 236868 397764
rect 236932 397762 236938 397764
rect 237189 397762 237255 397765
rect 236932 397760 237255 397762
rect 236932 397704 237194 397760
rect 237250 397704 237255 397760
rect 236932 397702 237255 397704
rect 236932 397700 236938 397702
rect 237189 397699 237255 397702
rect 237966 397700 237972 397764
rect 238036 397762 238042 397764
rect 238477 397762 238543 397765
rect 238036 397760 238543 397762
rect 238036 397704 238482 397760
rect 238538 397704 238543 397760
rect 238036 397702 238543 397704
rect 238036 397700 238042 397702
rect 238477 397699 238543 397702
rect 239673 397762 239739 397765
rect 239990 397762 239996 397764
rect 239673 397760 239996 397762
rect 239673 397704 239678 397760
rect 239734 397704 239996 397760
rect 239673 397702 239996 397704
rect 239673 397699 239739 397702
rect 239990 397700 239996 397702
rect 240060 397700 240066 397764
rect 242433 397762 242499 397765
rect 242750 397762 242756 397764
rect 242433 397760 242756 397762
rect 242433 397704 242438 397760
rect 242494 397704 242756 397760
rect 242433 397702 242756 397704
rect 242433 397699 242499 397702
rect 242750 397700 242756 397702
rect 242820 397700 242826 397764
rect 243670 397700 243676 397764
rect 243740 397762 243746 397764
rect 243997 397762 244063 397765
rect 243740 397760 244063 397762
rect 243740 397704 244002 397760
rect 244058 397704 244063 397760
rect 243740 397702 244063 397704
rect 243740 397700 243746 397702
rect 243997 397699 244063 397702
rect 246614 397700 246620 397764
rect 246684 397762 246690 397764
rect 246941 397762 247007 397765
rect 246684 397760 247007 397762
rect 246684 397704 246946 397760
rect 247002 397704 247007 397760
rect 246684 397702 247007 397704
rect 246684 397700 246690 397702
rect 246941 397699 247007 397702
rect 247718 397700 247724 397764
rect 247788 397762 247794 397764
rect 248137 397762 248203 397765
rect 247788 397760 248203 397762
rect 247788 397704 248142 397760
rect 248198 397704 248203 397760
rect 247788 397702 248203 397704
rect 247788 397700 247794 397702
rect 248137 397699 248203 397702
rect 248638 397700 248644 397764
rect 248708 397762 248714 397764
rect 249701 397762 249767 397765
rect 248708 397760 249767 397762
rect 248708 397704 249706 397760
rect 249762 397704 249767 397760
rect 248708 397702 249767 397704
rect 248708 397700 248714 397702
rect 249701 397699 249767 397702
rect 250478 397700 250484 397764
rect 250548 397762 250554 397764
rect 250989 397762 251055 397765
rect 250548 397760 251055 397762
rect 250548 397704 250994 397760
rect 251050 397704 251055 397760
rect 250548 397702 251055 397704
rect 250548 397700 250554 397702
rect 250989 397699 251055 397702
rect 251950 397700 251956 397764
rect 252020 397762 252026 397764
rect 252185 397762 252251 397765
rect 252020 397760 252251 397762
rect 252020 397704 252190 397760
rect 252246 397704 252251 397760
rect 252020 397702 252251 397704
rect 252020 397700 252026 397702
rect 252185 397699 252251 397702
rect 253238 397700 253244 397764
rect 253308 397762 253314 397764
rect 253749 397762 253815 397765
rect 253308 397760 253815 397762
rect 253308 397704 253754 397760
rect 253810 397704 253815 397760
rect 253308 397702 253815 397704
rect 253890 397762 253950 397838
rect 254710 397836 254716 397900
rect 254780 397898 254786 397900
rect 263542 397898 263548 397900
rect 254780 397838 263548 397898
rect 254780 397836 254786 397838
rect 263542 397836 263548 397838
rect 263612 397836 263618 397900
rect 261477 397762 261543 397765
rect 253890 397760 261543 397762
rect 253890 397704 261482 397760
rect 261538 397704 261543 397760
rect 253890 397702 261543 397704
rect 253308 397700 253314 397702
rect 253749 397699 253815 397702
rect 261477 397699 261543 397702
rect 214741 397624 215034 397626
rect 214741 397568 214746 397624
rect 214802 397568 215034 397624
rect 214741 397566 215034 397568
rect 215477 397628 215543 397629
rect 215477 397624 215524 397628
rect 215588 397626 215594 397628
rect 215477 397568 215482 397624
rect 214741 397563 214807 397566
rect 215477 397564 215524 397568
rect 215588 397566 215634 397626
rect 215588 397564 215594 397566
rect 216622 397564 216628 397628
rect 216692 397626 216698 397628
rect 216857 397626 216923 397629
rect 216692 397624 216923 397626
rect 216692 397568 216862 397624
rect 216918 397568 216923 397624
rect 216692 397566 216923 397568
rect 216692 397564 216698 397566
rect 215477 397563 215543 397564
rect 216857 397563 216923 397566
rect 218237 397626 218303 397629
rect 218830 397626 218836 397628
rect 218237 397624 218836 397626
rect 218237 397568 218242 397624
rect 218298 397568 218836 397624
rect 218237 397566 218836 397568
rect 218237 397563 218303 397566
rect 218830 397564 218836 397566
rect 218900 397564 218906 397628
rect 219525 397626 219591 397629
rect 219934 397626 219940 397628
rect 219525 397624 219940 397626
rect 219525 397568 219530 397624
rect 219586 397568 219940 397624
rect 219525 397566 219940 397568
rect 219525 397563 219591 397566
rect 219934 397564 219940 397566
rect 220004 397564 220010 397628
rect 220854 397564 220860 397628
rect 220924 397626 220930 397628
rect 221273 397626 221339 397629
rect 220924 397624 221339 397626
rect 220924 397568 221278 397624
rect 221334 397568 221339 397624
rect 220924 397566 221339 397568
rect 220924 397564 220930 397566
rect 221273 397563 221339 397566
rect 222377 397626 222443 397629
rect 223062 397626 223068 397628
rect 222377 397624 223068 397626
rect 222377 397568 222382 397624
rect 222438 397568 223068 397624
rect 222377 397566 223068 397568
rect 222377 397563 222443 397566
rect 223062 397564 223068 397566
rect 223132 397564 223138 397628
rect 223573 397626 223639 397629
rect 223798 397626 223804 397628
rect 223573 397624 223804 397626
rect 223573 397568 223578 397624
rect 223634 397568 223804 397624
rect 223573 397566 223804 397568
rect 223573 397563 223639 397566
rect 223798 397564 223804 397566
rect 223868 397564 223874 397628
rect 224953 397626 225019 397629
rect 225454 397626 225460 397628
rect 224953 397624 225460 397626
rect 224953 397568 224958 397624
rect 225014 397568 225460 397624
rect 224953 397566 225460 397568
rect 224953 397563 225019 397566
rect 225454 397564 225460 397566
rect 225524 397564 225530 397628
rect 228766 397564 228772 397628
rect 228836 397626 228842 397628
rect 229001 397626 229067 397629
rect 228836 397624 229067 397626
rect 228836 397568 229006 397624
rect 229062 397568 229067 397624
rect 228836 397566 229067 397568
rect 228836 397564 228842 397566
rect 229001 397563 229067 397566
rect 230054 397564 230060 397628
rect 230124 397626 230130 397628
rect 230381 397626 230447 397629
rect 230124 397624 230447 397626
rect 230124 397568 230386 397624
rect 230442 397568 230447 397624
rect 230124 397566 230447 397568
rect 230124 397564 230130 397566
rect 230381 397563 230447 397566
rect 230790 397564 230796 397628
rect 230860 397626 230866 397628
rect 231761 397626 231827 397629
rect 230860 397624 231827 397626
rect 230860 397568 231766 397624
rect 231822 397568 231827 397624
rect 230860 397566 231827 397568
rect 230860 397564 230866 397566
rect 231761 397563 231827 397566
rect 232814 397564 232820 397628
rect 232884 397626 232890 397628
rect 233141 397626 233207 397629
rect 232884 397624 233207 397626
rect 232884 397568 233146 397624
rect 233202 397568 233207 397624
rect 232884 397566 233207 397568
rect 232884 397564 232890 397566
rect 233141 397563 233207 397566
rect 234153 397626 234219 397629
rect 234286 397626 234292 397628
rect 234153 397624 234292 397626
rect 234153 397568 234158 397624
rect 234214 397568 234292 397624
rect 234153 397566 234292 397568
rect 234153 397563 234219 397566
rect 234286 397564 234292 397566
rect 234356 397564 234362 397628
rect 235390 397564 235396 397628
rect 235460 397626 235466 397628
rect 235717 397626 235783 397629
rect 235460 397624 235783 397626
rect 235460 397568 235722 397624
rect 235778 397568 235783 397624
rect 235460 397566 235783 397568
rect 235460 397564 235466 397566
rect 235717 397563 235783 397566
rect 237046 397564 237052 397628
rect 237116 397626 237122 397628
rect 237281 397626 237347 397629
rect 237116 397624 237347 397626
rect 237116 397568 237286 397624
rect 237342 397568 237347 397624
rect 237116 397566 237347 397568
rect 237116 397564 237122 397566
rect 237281 397563 237347 397566
rect 238150 397564 238156 397628
rect 238220 397626 238226 397628
rect 238385 397626 238451 397629
rect 238220 397624 238451 397626
rect 238220 397568 238390 397624
rect 238446 397568 238451 397624
rect 238220 397566 238451 397568
rect 238220 397564 238226 397566
rect 238385 397563 238451 397566
rect 239622 397564 239628 397628
rect 239692 397626 239698 397628
rect 239765 397626 239831 397629
rect 239692 397624 239831 397626
rect 239692 397568 239770 397624
rect 239826 397568 239831 397624
rect 239692 397566 239831 397568
rect 239692 397564 239698 397566
rect 239765 397563 239831 397566
rect 241094 397564 241100 397628
rect 241164 397626 241170 397628
rect 241421 397626 241487 397629
rect 241164 397624 241487 397626
rect 241164 397568 241426 397624
rect 241482 397568 241487 397624
rect 241164 397566 241487 397568
rect 241164 397564 241170 397566
rect 241421 397563 241487 397566
rect 242382 397564 242388 397628
rect 242452 397626 242458 397628
rect 242525 397626 242591 397629
rect 242452 397624 242591 397626
rect 242452 397568 242530 397624
rect 242586 397568 242591 397624
rect 242452 397566 242591 397568
rect 242452 397564 242458 397566
rect 242525 397563 242591 397566
rect 243854 397564 243860 397628
rect 243924 397626 243930 397628
rect 244181 397626 244247 397629
rect 243924 397624 244247 397626
rect 243924 397568 244186 397624
rect 244242 397568 244247 397624
rect 243924 397566 244247 397568
rect 243924 397564 243930 397566
rect 244181 397563 244247 397566
rect 244590 397564 244596 397628
rect 244660 397626 244666 397628
rect 245561 397626 245627 397629
rect 244660 397624 245627 397626
rect 244660 397568 245566 397624
rect 245622 397568 245627 397624
rect 244660 397566 245627 397568
rect 244660 397564 244666 397566
rect 245561 397563 245627 397566
rect 246430 397564 246436 397628
rect 246500 397626 246506 397628
rect 246665 397626 246731 397629
rect 246500 397624 246731 397626
rect 246500 397568 246670 397624
rect 246726 397568 246731 397624
rect 246500 397566 246731 397568
rect 246500 397564 246506 397566
rect 246665 397563 246731 397566
rect 248086 397564 248092 397628
rect 248156 397626 248162 397628
rect 248321 397626 248387 397629
rect 248156 397624 248387 397626
rect 248156 397568 248326 397624
rect 248382 397568 248387 397624
rect 248156 397566 248387 397568
rect 248156 397564 248162 397566
rect 248321 397563 248387 397566
rect 248822 397564 248828 397628
rect 248892 397626 248898 397628
rect 249517 397626 249583 397629
rect 248892 397624 249583 397626
rect 248892 397568 249522 397624
rect 249578 397568 249583 397624
rect 248892 397566 249583 397568
rect 248892 397564 248898 397566
rect 249517 397563 249583 397566
rect 250846 397564 250852 397628
rect 250916 397626 250922 397628
rect 251081 397626 251147 397629
rect 250916 397624 251147 397626
rect 250916 397568 251086 397624
rect 251142 397568 251147 397624
rect 250916 397566 251147 397568
rect 250916 397564 250922 397566
rect 251081 397563 251147 397566
rect 252134 397564 252140 397628
rect 252204 397626 252210 397628
rect 252277 397626 252343 397629
rect 252204 397624 252343 397626
rect 252204 397568 252282 397624
rect 252338 397568 252343 397624
rect 252204 397566 252343 397568
rect 252204 397564 252210 397566
rect 252277 397563 252343 397566
rect 253422 397564 253428 397628
rect 253492 397626 253498 397628
rect 253841 397626 253907 397629
rect 253492 397624 253907 397626
rect 253492 397568 253846 397624
rect 253902 397568 253907 397624
rect 253492 397566 253907 397568
rect 253492 397564 253498 397566
rect 253841 397563 253907 397566
rect 254710 397564 254716 397628
rect 254780 397626 254786 397628
rect 255129 397626 255195 397629
rect 254780 397624 255195 397626
rect 254780 397568 255134 397624
rect 255190 397568 255195 397624
rect 254780 397566 255195 397568
rect 254780 397564 254786 397566
rect 255129 397563 255195 397566
rect 211337 397492 211403 397493
rect 211286 397490 211292 397492
rect 206461 397488 210618 397490
rect 206461 397432 206466 397488
rect 206522 397432 210618 397488
rect 206461 397430 210618 397432
rect 211246 397430 211292 397490
rect 211356 397488 211403 397492
rect 212533 397492 212599 397493
rect 212717 397492 212783 397493
rect 214189 397492 214255 397493
rect 215385 397492 215451 397493
rect 215753 397492 215819 397493
rect 212533 397490 212580 397492
rect 211398 397432 211403 397488
rect 206461 397427 206527 397430
rect 211286 397428 211292 397430
rect 211356 397428 211403 397432
rect 212488 397488 212580 397490
rect 212488 397432 212538 397488
rect 212488 397430 212580 397432
rect 211337 397427 211403 397428
rect 212533 397428 212580 397430
rect 212644 397428 212650 397492
rect 212717 397488 212764 397492
rect 212828 397490 212834 397492
rect 212717 397432 212722 397488
rect 212717 397428 212764 397432
rect 212828 397430 212874 397490
rect 214189 397488 214236 397492
rect 214300 397490 214306 397492
rect 215334 397490 215340 397492
rect 214189 397432 214194 397488
rect 212828 397428 212834 397430
rect 214189 397428 214236 397432
rect 214300 397430 214346 397490
rect 215294 397430 215340 397490
rect 215404 397488 215451 397492
rect 215702 397490 215708 397492
rect 215446 397432 215451 397488
rect 214300 397428 214306 397430
rect 215334 397428 215340 397430
rect 215404 397428 215451 397432
rect 215662 397430 215708 397490
rect 215772 397488 215819 397492
rect 215814 397432 215819 397488
rect 215702 397428 215708 397430
rect 215772 397428 215819 397432
rect 216806 397428 216812 397492
rect 216876 397490 216882 397492
rect 216949 397490 217015 397493
rect 216876 397488 217015 397490
rect 216876 397432 216954 397488
rect 217010 397432 217015 397488
rect 216876 397430 217015 397432
rect 216876 397428 216882 397430
rect 212533 397427 212599 397428
rect 212717 397427 212783 397428
rect 214189 397427 214255 397428
rect 215385 397427 215451 397428
rect 215753 397427 215819 397428
rect 216949 397427 217015 397430
rect 218145 397490 218211 397493
rect 218646 397490 218652 397492
rect 218145 397488 218652 397490
rect 218145 397432 218150 397488
rect 218206 397432 218652 397488
rect 218145 397430 218652 397432
rect 218145 397427 218211 397430
rect 218646 397428 218652 397430
rect 218716 397428 218722 397492
rect 219566 397428 219572 397492
rect 219636 397490 219642 397492
rect 219893 397490 219959 397493
rect 219636 397488 219959 397490
rect 219636 397432 219898 397488
rect 219954 397432 219959 397488
rect 219636 397430 219959 397432
rect 219636 397428 219642 397430
rect 219893 397427 219959 397430
rect 220997 397492 221063 397493
rect 220997 397488 221044 397492
rect 221108 397490 221114 397492
rect 220997 397432 221002 397488
rect 220997 397428 221044 397432
rect 221108 397430 221154 397490
rect 221108 397428 221114 397430
rect 222142 397428 222148 397492
rect 222212 397490 222218 397492
rect 222285 397490 222351 397493
rect 222212 397488 222351 397490
rect 222212 397432 222290 397488
rect 222346 397432 222351 397488
rect 222212 397430 222351 397432
rect 222212 397428 222218 397430
rect 220997 397427 221063 397428
rect 222285 397427 222351 397430
rect 223849 397490 223915 397493
rect 223982 397490 223988 397492
rect 223849 397488 223988 397490
rect 223849 397432 223854 397488
rect 223910 397432 223988 397488
rect 223849 397430 223988 397432
rect 223849 397427 223915 397430
rect 223982 397428 223988 397430
rect 224052 397428 224058 397492
rect 225086 397428 225092 397492
rect 225156 397490 225162 397492
rect 225413 397490 225479 397493
rect 225156 397488 225479 397490
rect 225156 397432 225418 397488
rect 225474 397432 225479 397488
rect 225156 397430 225479 397432
rect 225156 397428 225162 397430
rect 225413 397427 225479 397430
rect 226374 397428 226380 397492
rect 226444 397490 226450 397492
rect 226517 397490 226583 397493
rect 226444 397488 226583 397490
rect 226444 397432 226522 397488
rect 226578 397432 226583 397488
rect 226444 397430 226583 397432
rect 226444 397428 226450 397430
rect 226517 397427 226583 397430
rect 228398 397428 228404 397492
rect 228468 397490 228474 397492
rect 228725 397490 228791 397493
rect 228909 397492 228975 397493
rect 228909 397490 228956 397492
rect 228468 397488 228791 397490
rect 228468 397432 228730 397488
rect 228786 397432 228791 397488
rect 228468 397430 228791 397432
rect 228864 397488 228956 397490
rect 228864 397432 228914 397488
rect 228864 397430 228956 397432
rect 228468 397428 228474 397430
rect 228725 397427 228791 397430
rect 228909 397428 228956 397430
rect 229020 397428 229026 397492
rect 230105 397490 230171 397493
rect 230238 397490 230244 397492
rect 230105 397488 230244 397490
rect 230105 397432 230110 397488
rect 230166 397432 230244 397488
rect 230105 397430 230244 397432
rect 228909 397427 228975 397428
rect 230105 397427 230171 397430
rect 230238 397428 230244 397430
rect 230308 397428 230314 397492
rect 230974 397428 230980 397492
rect 231044 397490 231050 397492
rect 231485 397490 231551 397493
rect 233049 397492 233115 397493
rect 232998 397490 233004 397492
rect 231044 397488 231551 397490
rect 231044 397432 231490 397488
rect 231546 397432 231551 397488
rect 231044 397430 231551 397432
rect 232958 397430 233004 397490
rect 233068 397488 233115 397492
rect 234061 397492 234127 397493
rect 234061 397490 234108 397492
rect 233110 397432 233115 397488
rect 231044 397428 231050 397430
rect 231485 397427 231551 397430
rect 232998 397428 233004 397430
rect 233068 397428 233115 397432
rect 234016 397488 234108 397490
rect 234016 397432 234066 397488
rect 234016 397430 234108 397432
rect 233049 397427 233115 397428
rect 234061 397428 234108 397430
rect 234172 397428 234178 397492
rect 234521 397490 234587 397493
rect 234521 397488 234630 397490
rect 234521 397432 234526 397488
rect 234582 397432 234630 397488
rect 234061 397427 234127 397428
rect 234521 397427 234630 397432
rect 235574 397428 235580 397492
rect 235644 397490 235650 397492
rect 235809 397490 235875 397493
rect 235644 397488 235875 397490
rect 235644 397432 235814 397488
rect 235870 397432 235875 397488
rect 235644 397430 235875 397432
rect 235644 397428 235650 397430
rect 235809 397427 235875 397430
rect 237097 397490 237163 397493
rect 237230 397490 237236 397492
rect 237097 397488 237236 397490
rect 237097 397432 237102 397488
rect 237158 397432 237236 397488
rect 237097 397430 237236 397432
rect 237097 397427 237163 397430
rect 237230 397428 237236 397430
rect 237300 397428 237306 397492
rect 238334 397428 238340 397492
rect 238404 397490 238410 397492
rect 238569 397490 238635 397493
rect 238404 397488 238635 397490
rect 238404 397432 238574 397488
rect 238630 397432 238635 397488
rect 238404 397430 238635 397432
rect 238404 397428 238410 397430
rect 238569 397427 238635 397430
rect 239806 397428 239812 397492
rect 239876 397490 239882 397492
rect 239949 397490 240015 397493
rect 241329 397492 241395 397493
rect 241278 397490 241284 397492
rect 239876 397488 240015 397490
rect 239876 397432 239954 397488
rect 240010 397432 240015 397488
rect 239876 397430 240015 397432
rect 241238 397430 241284 397490
rect 241348 397488 241395 397492
rect 241390 397432 241395 397488
rect 239876 397428 239882 397430
rect 239949 397427 240015 397430
rect 241278 397428 241284 397430
rect 241348 397428 241395 397432
rect 242566 397428 242572 397492
rect 242636 397490 242642 397492
rect 242709 397490 242775 397493
rect 244089 397492 244155 397493
rect 244038 397490 244044 397492
rect 242636 397488 242775 397490
rect 242636 397432 242714 397488
rect 242770 397432 242775 397488
rect 242636 397430 242775 397432
rect 243998 397430 244044 397490
rect 244108 397488 244155 397492
rect 245469 397492 245535 397493
rect 245469 397490 245516 397492
rect 244150 397432 244155 397488
rect 242636 397428 242642 397430
rect 241329 397427 241395 397428
rect 242709 397427 242775 397430
rect 244038 397428 244044 397430
rect 244108 397428 244155 397432
rect 245424 397488 245516 397490
rect 245424 397432 245474 397488
rect 245424 397430 245516 397432
rect 244089 397427 244155 397428
rect 245469 397428 245516 397430
rect 245580 397428 245586 397492
rect 246246 397428 246252 397492
rect 246316 397490 246322 397492
rect 246481 397490 246547 397493
rect 246849 397492 246915 397493
rect 246798 397490 246804 397492
rect 246316 397488 246547 397490
rect 246316 397432 246486 397488
rect 246542 397432 246547 397488
rect 246316 397430 246547 397432
rect 246758 397430 246804 397490
rect 246868 397488 246915 397492
rect 246910 397432 246915 397488
rect 246316 397428 246322 397430
rect 245469 397427 245535 397428
rect 246481 397427 246547 397430
rect 246798 397428 246804 397430
rect 246868 397428 246915 397432
rect 247902 397428 247908 397492
rect 247972 397490 247978 397492
rect 248045 397490 248111 397493
rect 248229 397492 248295 397493
rect 248229 397490 248276 397492
rect 247972 397488 248111 397490
rect 247972 397432 248050 397488
rect 248106 397432 248111 397488
rect 247972 397430 248111 397432
rect 248184 397488 248276 397490
rect 248184 397432 248234 397488
rect 248184 397430 248276 397432
rect 247972 397428 247978 397430
rect 246849 397427 246915 397428
rect 248045 397427 248111 397430
rect 248229 397428 248276 397430
rect 248340 397428 248346 397492
rect 249006 397428 249012 397492
rect 249076 397490 249082 397492
rect 249609 397490 249675 397493
rect 249076 397488 249675 397490
rect 249076 397432 249614 397488
rect 249670 397432 249675 397488
rect 249076 397430 249675 397432
rect 249076 397428 249082 397430
rect 248229 397427 248295 397428
rect 249609 397427 249675 397430
rect 250662 397428 250668 397492
rect 250732 397490 250738 397492
rect 250805 397490 250871 397493
rect 252369 397492 252435 397493
rect 252318 397490 252324 397492
rect 250732 397488 250871 397490
rect 250732 397432 250810 397488
rect 250866 397432 250871 397488
rect 250732 397430 250871 397432
rect 252278 397430 252324 397490
rect 252388 397488 252435 397492
rect 253565 397492 253631 397493
rect 253565 397490 253612 397492
rect 252430 397432 252435 397488
rect 250732 397428 250738 397430
rect 250805 397427 250871 397430
rect 252318 397428 252324 397430
rect 252388 397428 252435 397432
rect 253520 397488 253612 397490
rect 253520 397432 253570 397488
rect 253520 397430 253612 397432
rect 252369 397427 252435 397428
rect 253565 397428 253612 397430
rect 253676 397428 253682 397492
rect 254894 397428 254900 397492
rect 254964 397490 254970 397492
rect 255037 397490 255103 397493
rect 254964 397488 255103 397490
rect 254964 397432 255042 397488
rect 255098 397432 255103 397488
rect 254964 397430 255103 397432
rect 254964 397428 254970 397430
rect 253565 397427 253631 397428
rect 255037 397427 255103 397430
rect 234570 397354 234630 397427
rect 310513 397354 310579 397357
rect 234570 397352 310579 397354
rect 234570 397296 310518 397352
rect 310574 397296 310579 397352
rect 234570 397294 310579 397296
rect 310513 397291 310579 397294
rect 235625 397218 235691 397221
rect 324313 397218 324379 397221
rect 235625 397216 324379 397218
rect 235625 397160 235630 397216
rect 235686 397160 324318 397216
rect 324374 397160 324379 397216
rect 235625 397158 324379 397160
rect 235625 397155 235691 397158
rect 324313 397155 324379 397158
rect 205633 397082 205699 397085
rect 226333 397082 226399 397085
rect 205633 397080 226399 397082
rect 205633 397024 205638 397080
rect 205694 397024 226338 397080
rect 226394 397024 226399 397080
rect 205633 397022 226399 397024
rect 205633 397019 205699 397022
rect 226333 397019 226399 397022
rect 235901 397082 235967 397085
rect 328453 397082 328519 397085
rect 235901 397080 328519 397082
rect 235901 397024 235906 397080
rect 235962 397024 328458 397080
rect 328514 397024 328519 397080
rect 235901 397022 328519 397024
rect 235901 397019 235967 397022
rect 328453 397019 328519 397022
rect 191833 396946 191899 396949
rect 225229 396946 225295 396949
rect 191833 396944 225295 396946
rect 191833 396888 191838 396944
rect 191894 396888 225234 396944
rect 225290 396888 225295 396944
rect 191833 396886 225295 396888
rect 191833 396883 191899 396886
rect 225229 396883 225295 396886
rect 238661 396946 238727 396949
rect 364333 396946 364399 396949
rect 238661 396944 364399 396946
rect 238661 396888 238666 396944
rect 238722 396888 364338 396944
rect 364394 396888 364399 396944
rect 238661 396886 364399 396888
rect 238661 396883 238727 396886
rect 364333 396883 364399 396886
rect 138013 396810 138079 396813
rect 221089 396810 221155 396813
rect 138013 396808 221155 396810
rect 138013 396752 138018 396808
rect 138074 396752 221094 396808
rect 221150 396752 221155 396808
rect 138013 396750 221155 396752
rect 138013 396747 138079 396750
rect 221089 396747 221155 396750
rect 242617 396810 242683 396813
rect 416773 396810 416839 396813
rect 242617 396808 416839 396810
rect 242617 396752 242622 396808
rect 242678 396752 416778 396808
rect 416834 396752 416839 396808
rect 242617 396750 416839 396752
rect 242617 396747 242683 396750
rect 416773 396747 416839 396750
rect 48313 396674 48379 396677
rect 214005 396674 214071 396677
rect 48313 396672 214071 396674
rect 48313 396616 48318 396672
rect 48374 396616 214010 396672
rect 214066 396616 214071 396672
rect 48313 396614 214071 396616
rect 48313 396611 48379 396614
rect 214005 396611 214071 396614
rect 255262 396612 255268 396676
rect 255332 396674 255338 396676
rect 576853 396674 576919 396677
rect 255332 396672 576919 396674
rect 255332 396616 576858 396672
rect 576914 396616 576919 396672
rect 255332 396614 576919 396616
rect 255332 396612 255338 396614
rect 576853 396611 576919 396614
rect 232865 396538 232931 396541
rect 289813 396538 289879 396541
rect 232865 396536 289879 396538
rect 232865 396480 232870 396536
rect 232926 396480 289818 396536
rect 289874 396480 289879 396536
rect 232865 396478 289879 396480
rect 232865 396475 232931 396478
rect 289813 396475 289879 396478
rect 121453 395858 121519 395861
rect 219341 395858 219407 395861
rect 121453 395856 219407 395858
rect 121453 395800 121458 395856
rect 121514 395800 219346 395856
rect 219402 395800 219407 395856
rect 121453 395798 219407 395800
rect 121453 395795 121519 395798
rect 219341 395795 219407 395798
rect 118693 395722 118759 395725
rect 219750 395722 219756 395724
rect 118693 395720 219756 395722
rect 118693 395664 118698 395720
rect 118754 395664 219756 395720
rect 118693 395662 219756 395664
rect 118693 395659 118759 395662
rect 219750 395660 219756 395662
rect 219820 395660 219826 395724
rect 230422 395660 230428 395724
rect 230492 395722 230498 395724
rect 255589 395722 255655 395725
rect 230492 395720 255655 395722
rect 230492 395664 255594 395720
rect 255650 395664 255655 395720
rect 230492 395662 255655 395664
rect 230492 395660 230498 395662
rect 255589 395659 255655 395662
rect 67633 395586 67699 395589
rect 215886 395586 215892 395588
rect 67633 395584 215892 395586
rect 67633 395528 67638 395584
rect 67694 395528 215892 395584
rect 67633 395526 215892 395528
rect 67633 395523 67699 395526
rect 215886 395524 215892 395526
rect 215956 395524 215962 395588
rect 231577 395586 231643 395589
rect 273253 395586 273319 395589
rect 231577 395584 273319 395586
rect 231577 395528 231582 395584
rect 231638 395528 273258 395584
rect 273314 395528 273319 395584
rect 231577 395526 273319 395528
rect 231577 395523 231643 395526
rect 273253 395523 273319 395526
rect 27613 395450 27679 395453
rect 212574 395450 212580 395452
rect 27613 395448 212580 395450
rect 27613 395392 27618 395448
rect 27674 395392 212580 395448
rect 27613 395390 212580 395392
rect 27613 395387 27679 395390
rect 212574 395388 212580 395390
rect 212644 395388 212650 395452
rect 251030 395388 251036 395452
rect 251100 395450 251106 395452
rect 521653 395450 521719 395453
rect 251100 395448 521719 395450
rect 251100 395392 521658 395448
rect 521714 395392 521719 395448
rect 251100 395390 521719 395392
rect 251100 395388 251106 395390
rect 521653 395387 521719 395390
rect 11053 395314 11119 395317
rect 211153 395314 211219 395317
rect 11053 395312 211219 395314
rect 11053 395256 11058 395312
rect 11114 395256 211158 395312
rect 211214 395256 211219 395312
rect 11053 395254 211219 395256
rect 11053 395251 11119 395254
rect 211153 395251 211219 395254
rect 253054 395252 253060 395316
rect 253124 395314 253130 395316
rect 556153 395314 556219 395317
rect 253124 395312 556219 395314
rect 253124 395256 556158 395312
rect 556214 395256 556219 395312
rect 253124 395254 556219 395256
rect 253124 395252 253130 395254
rect 556153 395251 556219 395254
rect 208393 394362 208459 394365
rect 226374 394362 226380 394364
rect 208393 394360 226380 394362
rect 208393 394304 208398 394360
rect 208454 394304 226380 394360
rect 208393 394302 226380 394304
rect 208393 394299 208459 394302
rect 226374 394300 226380 394302
rect 226444 394300 226450 394364
rect 154573 394226 154639 394229
rect 223062 394226 223068 394228
rect 154573 394224 223068 394226
rect 154573 394168 154578 394224
rect 154634 394168 223068 394224
rect 154573 394166 223068 394168
rect 154573 394163 154639 394166
rect 223062 394164 223068 394166
rect 223132 394164 223138 394228
rect 82813 394090 82879 394093
rect 217174 394090 217180 394092
rect 82813 394088 217180 394090
rect 82813 394032 82818 394088
rect 82874 394032 217180 394088
rect 82813 394030 217180 394032
rect 82813 394027 82879 394030
rect 217174 394028 217180 394030
rect 217244 394028 217250 394092
rect 232129 394090 232195 394093
rect 232129 394088 232330 394090
rect 232129 394032 232134 394088
rect 232190 394032 232330 394088
rect 232129 394030 232330 394032
rect 232129 394027 232195 394030
rect 46933 393954 46999 393957
rect 214414 393954 214420 393956
rect 46933 393952 214420 393954
rect 46933 393896 46938 393952
rect 46994 393896 214420 393952
rect 46933 393894 214420 393896
rect 46933 393891 46999 393894
rect 214414 393892 214420 393894
rect 214484 393892 214490 393956
rect 232270 393821 232330 394030
rect 235390 393892 235396 393956
rect 235460 393954 235466 393956
rect 325693 393954 325759 393957
rect 235460 393952 325759 393954
rect 235460 393896 325698 393952
rect 325754 393896 325759 393952
rect 235460 393894 325759 393896
rect 235460 393892 235466 393894
rect 325693 393891 325759 393894
rect 232270 393816 232379 393821
rect 232270 393760 232318 393816
rect 232374 393760 232379 393816
rect 232270 393758 232379 393760
rect 232313 393755 232379 393758
rect 234889 393818 234955 393821
rect 235257 393818 235323 393821
rect 234889 393816 235323 393818
rect 234889 393760 234894 393816
rect 234950 393760 235262 393816
rect 235318 393760 235323 393816
rect 234889 393758 235323 393760
rect 234889 393755 234955 393758
rect 235257 393755 235323 393758
rect 583520 391628 584960 391868
rect 233509 389602 233575 389605
rect 233374 389600 233575 389602
rect 233374 389544 233514 389600
rect 233570 389544 233575 389600
rect 233374 389542 233575 389544
rect 233374 389197 233434 389542
rect 233509 389539 233575 389542
rect 233374 389192 233483 389197
rect 233374 389136 233422 389192
rect 233478 389136 233483 389192
rect 233374 389134 233483 389136
rect 233417 389131 233483 389134
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 236862 355540 236868 355604
rect 236932 355602 236938 355604
rect 345013 355602 345079 355605
rect 236932 355600 345079 355602
rect 236932 355544 345018 355600
rect 345074 355544 345079 355600
rect 236932 355542 345079 355544
rect 236932 355540 236938 355542
rect 345013 355539 345079 355542
rect 238150 355404 238156 355468
rect 238220 355466 238226 355468
rect 360193 355466 360259 355469
rect 238220 355464 360259 355466
rect 238220 355408 360198 355464
rect 360254 355408 360259 355464
rect 238220 355406 360259 355408
rect 238220 355404 238226 355406
rect 360193 355403 360259 355406
rect 30373 355330 30439 355333
rect 212758 355330 212764 355332
rect 30373 355328 212764 355330
rect 30373 355272 30378 355328
rect 30434 355272 212764 355328
rect 30373 355270 212764 355272
rect 30373 355267 30439 355270
rect 212758 355268 212764 355270
rect 212828 355268 212834 355332
rect 248638 355268 248644 355332
rect 248708 355330 248714 355332
rect 506473 355330 506539 355333
rect 248708 355328 506539 355330
rect 248708 355272 506478 355328
rect 506534 355272 506539 355328
rect 248708 355270 506539 355272
rect 248708 355268 248714 355270
rect 506473 355267 506539 355270
rect 234102 354316 234108 354380
rect 234172 354378 234178 354380
rect 304993 354378 305059 354381
rect 234172 354376 305059 354378
rect 234172 354320 304998 354376
rect 305054 354320 305059 354376
rect 234172 354318 305059 354320
rect 234172 354316 234178 354318
rect 304993 354315 305059 354318
rect 156597 354242 156663 354245
rect 219014 354242 219020 354244
rect 156597 354240 219020 354242
rect 156597 354184 156602 354240
rect 156658 354184 219020 354240
rect 156597 354182 219020 354184
rect 156597 354179 156663 354182
rect 219014 354180 219020 354182
rect 219084 354180 219090 354244
rect 243486 354180 243492 354244
rect 243556 354242 243562 354244
rect 431953 354242 432019 354245
rect 243556 354240 432019 354242
rect 243556 354184 431958 354240
rect 432014 354184 432019 354240
rect 243556 354182 432019 354184
rect 243556 354180 243562 354182
rect 431953 354179 432019 354182
rect 127617 354106 127683 354109
rect 215702 354106 215708 354108
rect 127617 354104 215708 354106
rect 127617 354048 127622 354104
rect 127678 354048 215708 354104
rect 127617 354046 215708 354048
rect 127617 354043 127683 354046
rect 215702 354044 215708 354046
rect 215772 354044 215778 354108
rect 244590 354044 244596 354108
rect 244660 354106 244666 354108
rect 452653 354106 452719 354109
rect 244660 354104 452719 354106
rect 244660 354048 452658 354104
rect 452714 354048 452719 354104
rect 244660 354046 452719 354048
rect 244660 354044 244666 354046
rect 452653 354043 452719 354046
rect 11145 353970 11211 353973
rect 211470 353970 211476 353972
rect 11145 353968 211476 353970
rect 11145 353912 11150 353968
rect 11206 353912 211476 353968
rect 11145 353910 211476 353912
rect 11145 353907 11211 353910
rect 211470 353908 211476 353910
rect 211540 353908 211546 353972
rect 228582 353908 228588 353972
rect 228652 353970 228658 353972
rect 237925 353970 237991 353973
rect 228652 353968 237991 353970
rect 228652 353912 237930 353968
rect 237986 353912 237991 353968
rect 228652 353910 237991 353912
rect 228652 353908 228658 353910
rect 237925 353907 237991 353910
rect 253238 353908 253244 353972
rect 253308 353970 253314 353972
rect 557533 353970 557599 353973
rect 253308 353968 557599 353970
rect 253308 353912 557538 353968
rect 557594 353912 557599 353968
rect 253308 353910 557599 353912
rect 253308 353908 253314 353910
rect 557533 353907 557599 353910
rect 229870 353500 229876 353564
rect 229940 353562 229946 353564
rect 236637 353562 236703 353565
rect 229940 353560 236703 353562
rect 229940 353504 236642 353560
rect 236698 353504 236703 353560
rect 229940 353502 236703 353504
rect 229940 353500 229946 353502
rect 236637 353499 236703 353502
rect 228398 353364 228404 353428
rect 228468 353426 228474 353428
rect 231117 353426 231183 353429
rect 228468 353424 231183 353426
rect 228468 353368 231122 353424
rect 231178 353368 231183 353424
rect 228468 353366 231183 353368
rect 228468 353364 228474 353366
rect 231117 353363 231183 353366
rect 187693 353018 187759 353021
rect 225086 353018 225092 353020
rect 187693 353016 225092 353018
rect 187693 352960 187698 353016
rect 187754 352960 225092 353016
rect 187693 352958 225092 352960
rect 187693 352955 187759 352958
rect 225086 352956 225092 352958
rect 225156 352956 225162 353020
rect 237046 352956 237052 353020
rect 237116 353018 237122 353020
rect 346393 353018 346459 353021
rect 237116 353016 346459 353018
rect 237116 352960 346398 353016
rect 346454 352960 346459 353016
rect 237116 352958 346459 352960
rect 237116 352956 237122 352958
rect 346393 352955 346459 352958
rect 172513 352882 172579 352885
rect 224166 352882 224172 352884
rect 172513 352880 224172 352882
rect 172513 352824 172518 352880
rect 172574 352824 224172 352880
rect 172513 352822 224172 352824
rect 172513 352819 172579 352822
rect 224166 352820 224172 352822
rect 224236 352820 224242 352884
rect 242382 352820 242388 352884
rect 242452 352882 242458 352884
rect 414013 352882 414079 352885
rect 242452 352880 414079 352882
rect 242452 352824 414018 352880
rect 414074 352824 414079 352880
rect 242452 352822 414079 352824
rect 242452 352820 242458 352822
rect 414013 352819 414079 352822
rect 135253 352746 135319 352749
rect 221222 352746 221228 352748
rect 135253 352744 221228 352746
rect 135253 352688 135258 352744
rect 135314 352688 221228 352744
rect 135253 352686 221228 352688
rect 135253 352683 135319 352686
rect 221222 352684 221228 352686
rect 221292 352684 221298 352748
rect 247718 352684 247724 352748
rect 247788 352746 247794 352748
rect 485773 352746 485839 352749
rect 247788 352744 485839 352746
rect 247788 352688 485778 352744
rect 485834 352688 485839 352744
rect 247788 352686 485839 352688
rect 247788 352684 247794 352686
rect 485773 352683 485839 352686
rect 122833 352610 122899 352613
rect 219566 352610 219572 352612
rect 122833 352608 219572 352610
rect 122833 352552 122838 352608
rect 122894 352552 219572 352608
rect 122833 352550 219572 352552
rect 122833 352547 122899 352550
rect 219566 352548 219572 352550
rect 219636 352548 219642 352612
rect 251766 352548 251772 352612
rect 251836 352610 251842 352612
rect 540973 352610 541039 352613
rect 251836 352608 541039 352610
rect 251836 352552 540978 352608
rect 541034 352552 541039 352608
rect 251836 352550 541039 352552
rect 251836 352548 251842 352550
rect 540973 352547 541039 352550
rect 255814 351868 255820 351932
rect 255884 351930 255890 351932
rect 583520 351930 584960 352020
rect 255884 351870 584960 351930
rect 255884 351868 255890 351870
rect 583520 351780 584960 351870
rect 153193 351386 153259 351389
rect 222142 351386 222148 351388
rect 153193 351384 222148 351386
rect 153193 351328 153198 351384
rect 153254 351328 222148 351384
rect 153193 351326 222148 351328
rect 153193 351323 153259 351326
rect 222142 351324 222148 351326
rect 222212 351324 222218 351388
rect 118785 351250 118851 351253
rect 219934 351250 219940 351252
rect 118785 351248 219940 351250
rect 118785 351192 118790 351248
rect 118846 351192 219940 351248
rect 118785 351190 219940 351192
rect 118785 351187 118851 351190
rect 219934 351188 219940 351190
rect 220004 351188 220010 351252
rect 241094 351188 241100 351252
rect 241164 351250 241170 351252
rect 398833 351250 398899 351253
rect 241164 351248 398899 351250
rect 241164 351192 398838 351248
rect 398894 351192 398899 351248
rect 241164 351190 398899 351192
rect 241164 351188 241170 351190
rect 398833 351187 398899 351190
rect 49693 351114 49759 351117
rect 214230 351114 214236 351116
rect 49693 351112 214236 351114
rect 49693 351056 49698 351112
rect 49754 351056 214236 351112
rect 49693 351054 214236 351056
rect 49693 351051 49759 351054
rect 214230 351052 214236 351054
rect 214300 351052 214306 351116
rect 251950 351052 251956 351116
rect 252020 351114 252026 351116
rect 538213 351114 538279 351117
rect 252020 351112 538279 351114
rect 252020 351056 538218 351112
rect 538274 351056 538279 351112
rect 252020 351054 538279 351056
rect 252020 351052 252026 351054
rect 538213 351051 538279 351054
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 583520 298754 584960 298844
rect 583342 298694 584960 298754
rect 583342 298618 583402 298694
rect 583520 298618 584960 298694
rect 583342 298604 584960 298618
rect 583342 298558 583586 298604
rect 262622 298148 262628 298212
rect 262692 298210 262698 298212
rect 583526 298210 583586 298558
rect 262692 298150 583586 298210
rect 262692 298148 262698 298150
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3693 188866 3759 188869
rect -960 188864 3759 188866
rect -960 188808 3698 188864
rect 3754 188808 3759 188864
rect -960 188806 3759 188808
rect -960 188716 480 188806
rect 3693 188803 3759 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect 85573 177442 85639 177445
rect 216806 177442 216812 177444
rect 85573 177440 216812 177442
rect 85573 177384 85578 177440
rect 85634 177384 216812 177440
rect 85573 177382 216812 177384
rect 85573 177379 85639 177382
rect 216806 177380 216812 177382
rect 216876 177380 216882 177444
rect 81433 177306 81499 177309
rect 216990 177306 216996 177308
rect 81433 177304 216996 177306
rect 81433 177248 81438 177304
rect 81494 177248 216996 177304
rect 81433 177246 216996 177248
rect 81433 177243 81499 177246
rect 216990 177244 216996 177246
rect 217060 177244 217066 177308
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 232630 87620 232636 87684
rect 232700 87682 232706 87684
rect 291193 87682 291259 87685
rect 232700 87680 291259 87682
rect 232700 87624 291198 87680
rect 291254 87624 291259 87680
rect 232700 87622 291259 87624
rect 232700 87620 232706 87622
rect 291193 87619 291259 87622
rect 243670 87484 243676 87548
rect 243740 87546 243746 87548
rect 432045 87546 432111 87549
rect 243740 87544 432111 87546
rect 243740 87488 432050 87544
rect 432106 87488 432111 87544
rect 243740 87486 432111 87488
rect 243740 87484 243746 87486
rect 432045 87483 432111 87486
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 260598 45596 260604 45660
rect 260668 45658 260674 45660
rect 583526 45658 583586 46142
rect 260668 45598 583586 45658
rect 260668 45596 260674 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 246246 26828 246252 26892
rect 246316 26890 246322 26892
rect 465073 26890 465139 26893
rect 246316 26888 465139 26890
rect 246316 26832 465078 26888
rect 465134 26832 465139 26888
rect 246316 26830 465139 26832
rect 246316 26828 246322 26830
rect 465073 26827 465139 26830
rect 237230 25468 237236 25532
rect 237300 25530 237306 25532
rect 343633 25530 343699 25533
rect 237300 25528 343699 25530
rect 237300 25472 343638 25528
rect 343694 25472 343699 25528
rect 237300 25470 343699 25472
rect 237300 25468 237306 25470
rect 343633 25467 343699 25470
rect 252134 24244 252140 24308
rect 252204 24306 252210 24308
rect 539593 24306 539659 24309
rect 252204 24304 539659 24306
rect 252204 24248 539598 24304
rect 539654 24248 539659 24304
rect 252204 24246 539659 24248
rect 252204 24244 252210 24246
rect 539593 24243 539659 24246
rect 254894 24108 254900 24172
rect 254964 24170 254970 24172
rect 574093 24170 574159 24173
rect 254964 24168 574159 24170
rect 254964 24112 574098 24168
rect 574154 24112 574159 24168
rect 254964 24110 574159 24112
rect 254964 24108 254970 24110
rect 574093 24107 574159 24110
rect 246430 22748 246436 22812
rect 246500 22810 246506 22812
rect 466453 22810 466519 22813
rect 246500 22808 466519 22810
rect 246500 22752 466458 22808
rect 466514 22752 466519 22808
rect 246500 22750 466519 22752
rect 246500 22748 246506 22750
rect 466453 22747 466519 22750
rect 248822 22612 248828 22676
rect 248892 22674 248898 22676
rect 503713 22674 503779 22677
rect 248892 22672 503779 22674
rect 248892 22616 503718 22672
rect 503774 22616 503779 22672
rect 248892 22614 503779 22616
rect 248892 22612 248898 22614
rect 503713 22611 503779 22614
rect 243854 21252 243860 21316
rect 243924 21314 243930 21316
rect 434713 21314 434779 21317
rect 243924 21312 434779 21314
rect 243924 21256 434718 21312
rect 434774 21256 434779 21312
rect 243924 21254 434779 21256
rect 243924 21252 243930 21254
rect 434713 21251 434779 21254
rect 239622 20164 239628 20228
rect 239692 20226 239698 20228
rect 378133 20226 378199 20229
rect 239692 20224 378199 20226
rect 239692 20168 378138 20224
rect 378194 20168 378199 20224
rect 239692 20166 378199 20168
rect 239692 20164 239698 20166
rect 378133 20163 378199 20166
rect 239438 20028 239444 20092
rect 239508 20090 239514 20092
rect 382365 20090 382431 20093
rect 239508 20088 382431 20090
rect 239508 20032 382370 20088
rect 382426 20032 382431 20088
rect 239508 20030 382431 20032
rect 239508 20028 239514 20030
rect 382365 20027 382431 20030
rect 246614 19892 246620 19956
rect 246684 19954 246690 19956
rect 470593 19954 470659 19957
rect 246684 19952 470659 19954
rect 246684 19896 470598 19952
rect 470654 19896 470659 19952
rect 246684 19894 470659 19896
rect 246684 19892 246690 19894
rect 470593 19891 470659 19894
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 298502 19348 298508 19412
rect 298572 19410 298578 19412
rect 583526 19410 583586 19622
rect 298572 19350 583586 19410
rect 298572 19348 298578 19350
rect 232814 18532 232820 18596
rect 232884 18594 232890 18596
rect 292573 18594 292639 18597
rect 232884 18592 292639 18594
rect 232884 18536 292578 18592
rect 292634 18536 292639 18592
rect 232884 18534 292639 18536
rect 232884 18532 232890 18534
rect 292573 18531 292639 18534
rect 230790 17444 230796 17508
rect 230860 17506 230866 17508
rect 276105 17506 276171 17509
rect 230860 17504 276171 17506
rect 230860 17448 276110 17504
rect 276166 17448 276171 17504
rect 230860 17446 276171 17448
rect 230860 17444 230866 17446
rect 276105 17443 276171 17446
rect 253606 17308 253612 17372
rect 253676 17370 253682 17372
rect 556245 17370 556311 17373
rect 253676 17368 556311 17370
rect 253676 17312 556250 17368
rect 556306 17312 556311 17368
rect 253676 17310 556311 17312
rect 253676 17308 253682 17310
rect 556245 17307 556311 17310
rect 253422 17172 253428 17236
rect 253492 17234 253498 17236
rect 558913 17234 558979 17237
rect 253492 17232 558979 17234
rect 253492 17176 558918 17232
rect 558974 17176 558979 17232
rect 253492 17174 558979 17176
rect 253492 17172 253498 17174
rect 558913 17171 558979 17174
rect 250662 15948 250668 16012
rect 250732 16010 250738 16012
rect 520273 16010 520339 16013
rect 250732 16008 520339 16010
rect 250732 15952 520278 16008
rect 520334 15952 520339 16008
rect 250732 15950 520339 15952
rect 250732 15948 250738 15950
rect 520273 15947 520339 15950
rect 250846 15812 250852 15876
rect 250916 15874 250922 15876
rect 523769 15874 523835 15877
rect 250916 15872 523835 15874
rect 250916 15816 523774 15872
rect 523830 15816 523835 15872
rect 250916 15814 523835 15816
rect 250916 15812 250922 15814
rect 523769 15811 523835 15814
rect 246798 14724 246804 14788
rect 246868 14786 246874 14788
rect 469857 14786 469923 14789
rect 246868 14784 469923 14786
rect 246868 14728 469862 14784
rect 469918 14728 469923 14784
rect 246868 14726 469923 14728
rect 246868 14724 246874 14726
rect 469857 14723 469923 14726
rect 247902 14588 247908 14652
rect 247972 14650 247978 14652
rect 484761 14650 484827 14653
rect 247972 14648 484827 14650
rect 247972 14592 484766 14648
rect 484822 14592 484827 14648
rect 247972 14590 484827 14592
rect 247972 14588 247978 14590
rect 484761 14587 484827 14590
rect 102225 14514 102291 14517
rect 218830 14514 218836 14516
rect 102225 14512 218836 14514
rect 102225 14456 102230 14512
rect 102286 14456 218836 14512
rect 102225 14454 218836 14456
rect 102225 14451 102291 14454
rect 218830 14452 218836 14454
rect 218900 14452 218906 14516
rect 248086 14452 248092 14516
rect 248156 14514 248162 14516
rect 488809 14514 488875 14517
rect 248156 14512 488875 14514
rect 248156 14456 488814 14512
rect 488870 14456 488875 14512
rect 248156 14454 488875 14456
rect 248156 14452 248162 14454
rect 488809 14451 488875 14454
rect 140037 13290 140103 13293
rect 216622 13290 216628 13292
rect 140037 13288 216628 13290
rect 140037 13232 140042 13288
rect 140098 13232 216628 13288
rect 140037 13230 216628 13232
rect 140037 13227 140103 13230
rect 216622 13228 216628 13230
rect 216692 13228 216698 13292
rect 66713 13154 66779 13157
rect 215518 13154 215524 13156
rect 66713 13152 215524 13154
rect 66713 13096 66718 13152
rect 66774 13096 215524 13152
rect 66713 13094 215524 13096
rect 66713 13091 66779 13094
rect 215518 13092 215524 13094
rect 215588 13092 215594 13156
rect 244038 13092 244044 13156
rect 244108 13154 244114 13156
rect 433977 13154 434043 13157
rect 244108 13152 434043 13154
rect 244108 13096 433982 13152
rect 434038 13096 434043 13152
rect 244108 13094 434043 13096
rect 244108 13092 244114 13094
rect 433977 13091 434043 13094
rect 13537 13018 13603 13021
rect 211286 13018 211292 13020
rect 13537 13016 211292 13018
rect 13537 12960 13542 13016
rect 13598 12960 211292 13016
rect 13537 12958 211292 12960
rect 13537 12955 13603 12958
rect 211286 12956 211292 12958
rect 211356 12956 211362 13020
rect 245510 12956 245516 13020
rect 245580 13018 245586 13020
rect 451641 13018 451707 13021
rect 245580 13016 451707 13018
rect 245580 12960 451646 13016
rect 451702 12960 451707 13016
rect 245580 12958 451707 12960
rect 245580 12956 245586 12958
rect 451641 12955 451707 12958
rect 241278 11868 241284 11932
rect 241348 11930 241354 11932
rect 398925 11930 398991 11933
rect 241348 11928 398991 11930
rect 241348 11872 398930 11928
rect 398986 11872 398991 11928
rect 241348 11870 398991 11872
rect 241348 11868 241354 11870
rect 398925 11867 398991 11870
rect 242750 11732 242756 11796
rect 242820 11794 242826 11796
rect 412633 11794 412699 11797
rect 242820 11792 412699 11794
rect 242820 11736 412638 11792
rect 412694 11736 412699 11792
rect 242820 11734 412699 11736
rect 242820 11732 242826 11734
rect 412633 11731 412699 11734
rect 17033 11658 17099 11661
rect 211102 11658 211108 11660
rect 17033 11656 211108 11658
rect 17033 11600 17038 11656
rect 17094 11600 211108 11656
rect 17033 11598 211108 11600
rect 17033 11595 17099 11598
rect 211102 11596 211108 11598
rect 211172 11596 211178 11660
rect 242566 11596 242572 11660
rect 242636 11658 242642 11660
rect 415485 11658 415551 11661
rect 242636 11656 415551 11658
rect 242636 11600 415490 11656
rect 415546 11600 415551 11656
rect 242636 11598 415551 11600
rect 242636 11596 242642 11598
rect 415485 11595 415551 11598
rect 238334 10508 238340 10572
rect 238404 10570 238410 10572
rect 363505 10570 363571 10573
rect 238404 10568 363571 10570
rect 238404 10512 363510 10568
rect 363566 10512 363571 10568
rect 238404 10510 363571 10512
rect 238404 10508 238410 10510
rect 363505 10507 363571 10510
rect 100753 10434 100819 10437
rect 218646 10434 218652 10436
rect 100753 10432 218652 10434
rect 100753 10376 100758 10432
rect 100814 10376 218652 10432
rect 100753 10374 218652 10376
rect 100753 10371 100819 10374
rect 218646 10372 218652 10374
rect 218716 10372 218722 10436
rect 239990 10372 239996 10436
rect 240060 10434 240066 10436
rect 377673 10434 377739 10437
rect 240060 10432 377739 10434
rect 240060 10376 377678 10432
rect 377734 10376 377739 10432
rect 240060 10374 377739 10376
rect 240060 10372 240066 10374
rect 377673 10371 377739 10374
rect 65057 10298 65123 10301
rect 215334 10298 215340 10300
rect 65057 10296 215340 10298
rect 65057 10240 65062 10296
rect 65118 10240 215340 10296
rect 65057 10238 215340 10240
rect 65057 10235 65123 10238
rect 215334 10236 215340 10238
rect 215404 10236 215410 10300
rect 239806 10236 239812 10300
rect 239876 10298 239882 10300
rect 381169 10298 381235 10301
rect 239876 10296 381235 10298
rect 239876 10240 381174 10296
rect 381230 10240 381235 10296
rect 239876 10238 381235 10240
rect 239876 10236 239882 10238
rect 381169 10235 381235 10238
rect 174261 9074 174327 9077
rect 223982 9074 223988 9076
rect 174261 9072 223988 9074
rect 174261 9016 174266 9072
rect 174322 9016 223988 9072
rect 174261 9014 223988 9016
rect 174261 9011 174327 9014
rect 223982 9012 223988 9014
rect 224052 9012 224058 9076
rect 230974 9012 230980 9076
rect 231044 9074 231050 9076
rect 272425 9074 272491 9077
rect 231044 9072 272491 9074
rect 231044 9016 272430 9072
rect 272486 9016 272491 9072
rect 231044 9014 272491 9016
rect 231044 9012 231050 9014
rect 272425 9011 272491 9014
rect 51349 8938 51415 8941
rect 214046 8938 214052 8940
rect 51349 8936 214052 8938
rect 51349 8880 51354 8936
rect 51410 8880 214052 8936
rect 51349 8878 214052 8880
rect 51349 8875 51415 8878
rect 214046 8876 214052 8878
rect 214116 8876 214122 8940
rect 235574 8876 235580 8940
rect 235644 8938 235650 8940
rect 327993 8938 328059 8941
rect 235644 8936 328059 8938
rect 235644 8880 327998 8936
rect 328054 8880 328059 8936
rect 235644 8878 328059 8880
rect 235644 8876 235650 8878
rect 327993 8875 328059 8878
rect 170765 7850 170831 7853
rect 223798 7850 223804 7852
rect 170765 7848 223804 7850
rect 170765 7792 170770 7848
rect 170826 7792 223804 7848
rect 170765 7790 223804 7792
rect 170765 7787 170831 7790
rect 223798 7788 223804 7790
rect 223868 7788 223874 7852
rect 232998 7788 233004 7852
rect 233068 7850 233074 7852
rect 292573 7850 292639 7853
rect 233068 7848 292639 7850
rect 233068 7792 292578 7848
rect 292634 7792 292639 7848
rect 233068 7790 292639 7792
rect 233068 7788 233074 7790
rect 292573 7787 292639 7790
rect 141233 7714 141299 7717
rect 220854 7714 220860 7716
rect 141233 7712 220860 7714
rect 141233 7656 141238 7712
rect 141294 7656 220860 7712
rect 141233 7654 220860 7656
rect 141233 7651 141299 7654
rect 220854 7652 220860 7654
rect 220924 7652 220930 7716
rect 234286 7652 234292 7716
rect 234356 7714 234362 7716
rect 306741 7714 306807 7717
rect 234356 7712 306807 7714
rect 234356 7656 306746 7712
rect 306802 7656 306807 7712
rect 234356 7654 306807 7656
rect 234356 7652 234362 7654
rect 306741 7651 306807 7654
rect 137645 7578 137711 7581
rect 221038 7578 221044 7580
rect 137645 7576 221044 7578
rect 137645 7520 137650 7576
rect 137706 7520 221044 7576
rect 137645 7518 221044 7520
rect 137645 7515 137711 7518
rect 221038 7516 221044 7518
rect 221108 7516 221114 7580
rect 233918 7516 233924 7580
rect 233988 7578 233994 7580
rect 310237 7578 310303 7581
rect 233988 7576 310303 7578
rect 233988 7520 310242 7576
rect 310298 7520 310303 7576
rect 233988 7518 310303 7520
rect 233988 7516 233994 7518
rect 310237 7515 310303 7518
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect 583520 6476 584960 6566
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 194409 6218 194475 6221
rect 224902 6218 224908 6220
rect 194409 6216 224908 6218
rect 194409 6160 194414 6216
rect 194470 6160 224908 6216
rect 194409 6158 224908 6160
rect 194409 6155 194475 6158
rect 224902 6156 224908 6158
rect 224972 6156 224978 6220
rect 254710 6156 254716 6220
rect 254780 6218 254786 6220
rect 576301 6218 576367 6221
rect 254780 6216 576367 6218
rect 254780 6160 576306 6216
rect 576362 6160 576367 6216
rect 254780 6158 576367 6160
rect 254780 6156 254786 6158
rect 576301 6155 576367 6158
rect 230238 5340 230244 5404
rect 230308 5402 230314 5404
rect 254669 5402 254735 5405
rect 230308 5400 254735 5402
rect 230308 5344 254674 5400
rect 254730 5344 254735 5400
rect 230308 5342 254735 5344
rect 230308 5340 230314 5342
rect 254669 5339 254735 5342
rect 230054 5204 230060 5268
rect 230124 5266 230130 5268
rect 258257 5266 258323 5269
rect 230124 5264 258323 5266
rect 230124 5208 258262 5264
rect 258318 5208 258323 5264
rect 230124 5206 258323 5208
rect 230124 5204 230130 5206
rect 258257 5203 258323 5206
rect 237966 5068 237972 5132
rect 238036 5130 238042 5132
rect 362309 5130 362375 5133
rect 238036 5128 362375 5130
rect 238036 5072 362314 5128
rect 362370 5072 362375 5128
rect 238036 5070 362375 5072
rect 238036 5068 238042 5070
rect 362309 5067 362375 5070
rect 249006 4932 249012 4996
rect 249076 4994 249082 4996
rect 505369 4994 505435 4997
rect 249076 4992 505435 4994
rect 249076 4936 505374 4992
rect 505430 4936 505435 4992
rect 249076 4934 505435 4936
rect 249076 4932 249082 4934
rect 505369 4931 505435 4934
rect 565 4858 631 4861
rect 209814 4858 209820 4860
rect 565 4856 209820 4858
rect 565 4800 570 4856
rect 626 4800 209820 4856
rect 565 4798 209820 4800
rect 565 4795 631 4798
rect 209814 4796 209820 4798
rect 209884 4796 209890 4860
rect 252318 4796 252324 4860
rect 252388 4858 252394 4860
rect 540789 4858 540855 4861
rect 252388 4856 540855 4858
rect 252388 4800 540794 4856
rect 540850 4800 540855 4856
rect 252388 4798 540855 4800
rect 252388 4796 252394 4798
rect 540789 4795 540855 4798
rect 226190 3708 226196 3772
rect 226260 3770 226266 3772
rect 299657 3770 299723 3773
rect 226260 3768 299723 3770
rect 226260 3712 299662 3768
rect 299718 3712 299723 3768
rect 226260 3710 299723 3712
rect 226260 3708 226266 3710
rect 299657 3707 299723 3710
rect 248270 3572 248276 3636
rect 248340 3634 248346 3636
rect 487613 3634 487679 3637
rect 248340 3632 487679 3634
rect 248340 3576 487618 3632
rect 487674 3576 487679 3632
rect 248340 3574 487679 3576
rect 248340 3572 248346 3574
rect 487613 3571 487679 3574
rect 228950 3436 228956 3500
rect 229020 3498 229026 3500
rect 239305 3498 239371 3501
rect 229020 3496 239371 3498
rect 229020 3440 239310 3496
rect 239366 3440 239371 3496
rect 229020 3438 239371 3440
rect 229020 3436 229026 3438
rect 239305 3435 239371 3438
rect 250478 3436 250484 3500
rect 250548 3498 250554 3500
rect 523033 3498 523099 3501
rect 250548 3496 523099 3498
rect 250548 3440 523038 3496
rect 523094 3440 523099 3496
rect 250548 3438 523099 3440
rect 250548 3436 250554 3438
rect 523033 3435 523099 3438
rect 175457 3362 175523 3365
rect 223614 3362 223620 3364
rect 175457 3360 223620 3362
rect 175457 3304 175462 3360
rect 175518 3304 223620 3360
rect 175457 3302 223620 3304
rect 175457 3299 175523 3302
rect 223614 3300 223620 3302
rect 223684 3300 223690 3364
rect 228766 3300 228772 3364
rect 228836 3362 228842 3364
rect 240501 3362 240567 3365
rect 228836 3360 240567 3362
rect 228836 3304 240506 3360
rect 240562 3304 240567 3360
rect 228836 3302 240567 3304
rect 228836 3300 228842 3302
rect 240501 3299 240567 3302
rect 262070 3300 262076 3364
rect 262140 3362 262146 3364
rect 579797 3362 579863 3365
rect 262140 3360 579863 3362
rect 262140 3304 579802 3360
rect 579858 3304 579863 3360
rect 262140 3302 579863 3304
rect 262140 3300 262146 3302
rect 579797 3299 579863 3302
<< via3 >>
rect 282132 699756 282196 699820
rect 102364 597484 102428 597548
rect 105308 597484 105372 597548
rect 106228 597484 106292 597548
rect 110460 597484 110524 597548
rect 115612 597484 115676 597548
rect 120580 597484 120644 597548
rect 125548 597484 125612 597548
rect 130516 597484 130580 597548
rect 135484 597484 135548 597548
rect 140636 597544 140700 597548
rect 140636 597488 140686 597544
rect 140686 597488 140700 597544
rect 140636 597484 140700 597488
rect 210004 597544 210068 597548
rect 210004 597488 210018 597544
rect 210018 597488 210068 597544
rect 210004 597484 210068 597488
rect 212396 597544 212460 597548
rect 212396 597488 212410 597544
rect 212410 597488 212460 597544
rect 212396 597484 212460 597488
rect 213500 597484 213564 597548
rect 214788 597544 214852 597548
rect 214788 597488 214838 597544
rect 214838 597488 214852 597544
rect 214788 597484 214852 597488
rect 215708 597484 215772 597548
rect 219204 597484 219268 597548
rect 225460 597544 225524 597548
rect 225460 597488 225510 597544
rect 225510 597488 225524 597544
rect 225460 597484 225524 597488
rect 230612 597544 230676 597548
rect 230612 597488 230662 597544
rect 230662 597488 230676 597544
rect 230612 597484 230676 597488
rect 235580 597484 235644 597548
rect 240548 597544 240612 597548
rect 240548 597488 240562 597544
rect 240562 597488 240612 597544
rect 240548 597484 240612 597488
rect 245516 597544 245580 597548
rect 245516 597488 245530 597544
rect 245530 597488 245580 597544
rect 245516 597484 245580 597488
rect 250484 597544 250548 597548
rect 250484 597488 250534 597544
rect 250534 597488 250548 597544
rect 250484 597484 250548 597488
rect 320036 597544 320100 597548
rect 320036 597488 320050 597544
rect 320050 597488 320100 597544
rect 320036 597484 320100 597488
rect 322244 597544 322308 597548
rect 322244 597488 322294 597544
rect 322294 597488 322308 597544
rect 322244 597484 322308 597488
rect 323348 597544 323412 597548
rect 323348 597488 323398 597544
rect 323398 597488 323412 597544
rect 323348 597484 323412 597488
rect 324820 597544 324884 597548
rect 324820 597488 324834 597544
rect 324834 597488 324884 597544
rect 324820 597484 324884 597488
rect 325740 597484 325804 597548
rect 330524 597484 330588 597548
rect 335124 597484 335188 597548
rect 340460 597544 340524 597548
rect 340460 597488 340510 597544
rect 340510 597488 340524 597544
rect 340460 597484 340524 597488
rect 345612 597544 345676 597548
rect 345612 597488 345662 597544
rect 345662 597488 345676 597544
rect 345612 597484 345676 597488
rect 350396 597544 350460 597548
rect 350396 597488 350446 597544
rect 350446 597488 350460 597544
rect 350396 597484 350460 597488
rect 354444 597484 354508 597548
rect 360516 597544 360580 597548
rect 360516 597488 360566 597544
rect 360566 597488 360580 597544
rect 360516 597484 360580 597488
rect 429884 597484 429948 597548
rect 435588 597484 435652 597548
rect 445524 597484 445588 597548
rect 460428 597484 460492 597548
rect 92980 597348 93044 597412
rect 98868 597348 98932 597412
rect 208900 597348 208964 597412
rect 315252 597348 315316 597412
rect 321140 597348 321204 597412
rect 430988 597348 431052 597412
rect 440372 597348 440436 597412
rect 455460 597408 455524 597412
rect 455460 597352 455474 597408
rect 455474 597352 455524 597408
rect 455460 597348 455524 597352
rect 465396 597348 465460 597412
rect 97764 597212 97828 597276
rect 207612 597272 207676 597276
rect 207612 597216 207662 597272
rect 207662 597216 207676 597272
rect 207612 597212 207676 597216
rect 318932 597212 318996 597276
rect 428964 597212 429028 597276
rect 433380 597272 433444 597276
rect 433380 597216 433394 597272
rect 433394 597216 433444 597272
rect 433380 597212 433444 597216
rect 450492 597212 450556 597276
rect 94268 597076 94332 597140
rect 103284 597076 103348 597140
rect 105676 597076 105740 597140
rect 106412 597076 106476 597140
rect 215340 597076 215404 597140
rect 99972 596940 100036 597004
rect 101076 596940 101140 597004
rect 211108 596940 211172 597004
rect 104756 596864 104820 596868
rect 317644 597076 317708 597140
rect 427676 597076 427740 597140
rect 434668 597136 434732 597140
rect 434668 597080 434718 597136
rect 434718 597080 434732 597136
rect 434668 597076 434732 597080
rect 321140 596940 321204 597004
rect 104756 596808 104806 596864
rect 104806 596808 104820 596864
rect 104756 596804 104820 596808
rect 325372 596804 325436 596868
rect 435220 596940 435284 597004
rect 470364 596940 470428 597004
rect 431724 596804 431788 596868
rect 205404 596532 205468 596596
rect 202828 596456 202892 596460
rect 202828 596400 202878 596456
rect 202878 596400 202892 596456
rect 202828 596396 202892 596400
rect 422892 596396 422956 596460
rect 95372 596260 95436 596324
rect 204300 596320 204364 596324
rect 204300 596264 204314 596320
rect 204314 596264 204364 596320
rect 204300 596260 204364 596264
rect 312860 596260 312924 596324
rect 314332 596260 314396 596324
rect 424180 596260 424244 596324
rect 425284 596260 425348 596324
rect 407804 523636 407868 523700
rect 407804 489772 407868 489836
rect 110460 489424 110524 489428
rect 110460 489368 110510 489424
rect 110510 489368 110524 489424
rect 110460 489364 110524 489368
rect 325372 489152 325436 489156
rect 325372 489096 325386 489152
rect 325386 489096 325436 489152
rect 325372 489092 325436 489096
rect 92980 488472 93044 488476
rect 92980 488416 92994 488472
rect 92994 488416 93044 488472
rect 92980 488412 93044 488416
rect 94268 488472 94332 488476
rect 94268 488416 94282 488472
rect 94282 488416 94332 488472
rect 94268 488412 94332 488416
rect 97764 488472 97828 488476
rect 97764 488416 97814 488472
rect 97814 488416 97828 488472
rect 97764 488412 97828 488416
rect 98868 488412 98932 488476
rect 99972 488472 100036 488476
rect 99972 488416 100022 488472
rect 100022 488416 100036 488472
rect 99972 488412 100036 488416
rect 101076 488472 101140 488476
rect 101076 488416 101126 488472
rect 101126 488416 101140 488472
rect 101076 488412 101140 488416
rect 102364 488472 102428 488476
rect 102364 488416 102414 488472
rect 102414 488416 102428 488472
rect 102364 488412 102428 488416
rect 104756 488472 104820 488476
rect 104756 488416 104806 488472
rect 104806 488416 104820 488472
rect 104756 488412 104820 488416
rect 105308 488472 105372 488476
rect 105308 488416 105358 488472
rect 105358 488416 105372 488472
rect 105308 488412 105372 488416
rect 105676 488472 105740 488476
rect 105676 488416 105726 488472
rect 105726 488416 105740 488472
rect 105676 488412 105740 488416
rect 115612 488472 115676 488476
rect 115612 488416 115662 488472
rect 115662 488416 115676 488472
rect 115612 488412 115676 488416
rect 120580 488472 120644 488476
rect 120580 488416 120630 488472
rect 120630 488416 120644 488472
rect 120580 488412 120644 488416
rect 125548 488472 125612 488476
rect 125548 488416 125598 488472
rect 125598 488416 125612 488472
rect 125548 488412 125612 488416
rect 130516 488412 130580 488476
rect 135484 488472 135548 488476
rect 135484 488416 135534 488472
rect 135534 488416 135548 488472
rect 135484 488412 135548 488416
rect 140636 488472 140700 488476
rect 140636 488416 140686 488472
rect 140686 488416 140700 488472
rect 140636 488412 140700 488416
rect 95372 488336 95436 488340
rect 205404 488412 205468 488476
rect 215340 488472 215404 488476
rect 215340 488416 215354 488472
rect 215354 488416 215404 488472
rect 215340 488412 215404 488416
rect 220492 488412 220556 488476
rect 225460 488412 225524 488476
rect 230428 488472 230492 488476
rect 230428 488416 230478 488472
rect 230478 488416 230492 488472
rect 230428 488412 230492 488416
rect 330524 488472 330588 488476
rect 330524 488416 330538 488472
rect 330538 488416 330588 488472
rect 330524 488412 330588 488416
rect 335492 488472 335556 488476
rect 335492 488416 335506 488472
rect 335506 488416 335556 488472
rect 335492 488412 335556 488416
rect 340644 488472 340708 488476
rect 340644 488416 340658 488472
rect 340658 488416 340708 488472
rect 340644 488412 340708 488416
rect 345612 488412 345676 488476
rect 350396 488472 350460 488476
rect 350396 488416 350410 488472
rect 350410 488416 350460 488472
rect 350396 488412 350460 488416
rect 355548 488412 355612 488476
rect 360516 488472 360580 488476
rect 360516 488416 360530 488472
rect 360530 488416 360580 488472
rect 360516 488412 360580 488416
rect 422892 488412 422956 488476
rect 424180 488412 424244 488476
rect 435220 488412 435284 488476
rect 440372 488412 440436 488476
rect 445524 488412 445588 488476
rect 450492 488412 450556 488476
rect 95372 488280 95386 488336
rect 95386 488280 95436 488336
rect 95372 488276 95436 488280
rect 314332 488276 314396 488340
rect 315436 488140 315500 488204
rect 425284 488276 425348 488340
rect 430988 488276 431052 488340
rect 465396 488276 465460 488340
rect 428964 488140 429028 488204
rect 429884 488140 429948 488204
rect 435588 488140 435652 488204
rect 203012 488004 203076 488068
rect 204300 488064 204364 488068
rect 204300 488008 204314 488064
rect 204314 488008 204364 488064
rect 204300 488004 204364 488008
rect 212212 488004 212276 488068
rect 455460 488064 455524 488068
rect 455460 488008 455474 488064
rect 455474 488008 455524 488064
rect 455460 488004 455524 488008
rect 470732 488004 470796 488068
rect 211108 487928 211172 487932
rect 211108 487872 211158 487928
rect 211158 487872 211172 487928
rect 211108 487868 211172 487872
rect 235580 487928 235644 487932
rect 235580 487872 235630 487928
rect 235630 487872 235644 487928
rect 235580 487868 235644 487872
rect 240548 487868 240612 487932
rect 318932 487928 318996 487932
rect 318932 487872 318946 487928
rect 318946 487872 318996 487928
rect 318932 487868 318996 487872
rect 460428 487868 460492 487932
rect 427676 487732 427740 487796
rect 432276 487596 432340 487660
rect 103284 487460 103348 487524
rect 210004 487520 210068 487524
rect 210004 487464 210054 487520
rect 210054 487464 210068 487520
rect 210004 487460 210068 487464
rect 213316 487460 213380 487524
rect 250484 487520 250548 487524
rect 250484 487464 250498 487520
rect 250498 487464 250548 487520
rect 250484 487460 250548 487464
rect 205404 487324 205468 487388
rect 245516 487384 245580 487388
rect 245516 487328 245566 487384
rect 245566 487328 245580 487384
rect 245516 487324 245580 487328
rect 323348 487324 323412 487388
rect 433380 487384 433444 487388
rect 433380 487328 433394 487384
rect 433394 487328 433444 487384
rect 433380 487324 433444 487328
rect 203012 487188 203076 487252
rect 204300 487188 204364 487252
rect 207612 487248 207676 487252
rect 207612 487192 207662 487248
rect 207662 487192 207676 487248
rect 207612 487188 207676 487192
rect 208900 487188 208964 487252
rect 214788 487188 214852 487252
rect 215708 487188 215772 487252
rect 312860 487188 312924 487252
rect 317644 487188 317708 487252
rect 320036 487248 320100 487252
rect 320036 487192 320086 487248
rect 320086 487192 320100 487248
rect 320036 487188 320100 487192
rect 321140 487188 321204 487252
rect 322244 487248 322308 487252
rect 322244 487192 322258 487248
rect 322258 487192 322308 487248
rect 322244 487188 322308 487192
rect 324820 487248 324884 487252
rect 324820 487192 324870 487248
rect 324870 487192 324884 487248
rect 324820 487188 324884 487192
rect 325740 487188 325804 487252
rect 434852 487188 434916 487252
rect 282132 476716 282196 476780
rect 257476 446796 257540 446860
rect 262628 446660 262692 446724
rect 254532 446116 254596 446180
rect 298508 446116 298572 446180
rect 257292 445708 257356 445772
rect 254900 445572 254964 445636
rect 260604 445572 260668 445636
rect 254716 445028 254780 445092
rect 260052 444348 260116 444412
rect 253796 444076 253860 444140
rect 212948 443804 213012 443868
rect 232268 443864 232332 443868
rect 232268 443808 232318 443864
rect 232318 443808 232332 443864
rect 232268 443804 232332 443808
rect 233188 443864 233252 443868
rect 233188 443808 233238 443864
rect 233238 443808 233252 443864
rect 233188 443804 233252 443808
rect 234844 443864 234908 443868
rect 234844 443808 234894 443864
rect 234894 443808 234908 443864
rect 234844 443804 234908 443808
rect 210372 443396 210436 443460
rect 214236 443532 214300 443596
rect 255820 443532 255884 443596
rect 256556 443592 256620 443596
rect 256556 443536 256606 443592
rect 256606 443536 256620 443592
rect 256556 443532 256620 443536
rect 259132 443396 259196 443460
rect 259316 443456 259380 443460
rect 259316 443400 259366 443456
rect 259366 443400 259380 443456
rect 259316 443396 259380 443400
rect 262076 443456 262140 443460
rect 262076 443400 262126 443456
rect 262126 443400 262140 443456
rect 262076 443396 262140 443400
rect 214236 443260 214300 443324
rect 214420 443260 214484 443324
rect 210372 442988 210436 443052
rect 214420 442988 214484 443052
rect 232268 442580 232332 442644
rect 233188 442444 233252 442508
rect 234844 442308 234908 442372
rect 212948 442172 213012 442236
rect 383332 402868 383396 402932
rect 259132 401508 259196 401572
rect 383332 401508 383396 401572
rect 256556 400148 256620 400212
rect 253060 399468 253124 399532
rect 253796 399468 253860 399532
rect 253244 399332 253308 399396
rect 255268 399256 255332 399260
rect 255268 399200 255282 399256
rect 255282 399200 255332 399256
rect 255268 399196 255332 399200
rect 217180 398788 217244 398852
rect 253244 398712 253308 398716
rect 254532 399060 254596 399124
rect 257476 399060 257540 399124
rect 254900 398924 254964 398988
rect 253244 398656 253258 398712
rect 253258 398656 253308 398712
rect 253244 398652 253308 398656
rect 260052 398516 260116 398580
rect 209820 397700 209884 397764
rect 214420 397836 214484 397900
rect 211108 397700 211172 397764
rect 211476 397564 211540 397628
rect 214052 397564 214116 397628
rect 257292 398380 257356 398444
rect 263548 398380 263612 398444
rect 259316 398244 259380 398308
rect 226196 397972 226260 398036
rect 224172 397836 224236 397900
rect 230428 397836 230492 397900
rect 239444 397836 239508 397900
rect 243492 397836 243556 397900
rect 251036 397836 251100 397900
rect 251772 397836 251836 397900
rect 215892 397700 215956 397764
rect 216996 397700 217060 397764
rect 219020 397700 219084 397764
rect 219756 397700 219820 397764
rect 221228 397700 221292 397764
rect 223620 397700 223684 397764
rect 228588 397700 228652 397764
rect 229876 397700 229940 397764
rect 232636 397700 232700 397764
rect 233924 397700 233988 397764
rect 236868 397700 236932 397764
rect 237972 397700 238036 397764
rect 239996 397700 240060 397764
rect 242756 397700 242820 397764
rect 243676 397700 243740 397764
rect 246620 397700 246684 397764
rect 247724 397700 247788 397764
rect 248644 397700 248708 397764
rect 250484 397700 250548 397764
rect 251956 397700 252020 397764
rect 253244 397700 253308 397764
rect 254716 397836 254780 397900
rect 263548 397836 263612 397900
rect 215524 397624 215588 397628
rect 215524 397568 215538 397624
rect 215538 397568 215588 397624
rect 215524 397564 215588 397568
rect 216628 397564 216692 397628
rect 218836 397564 218900 397628
rect 219940 397564 220004 397628
rect 220860 397564 220924 397628
rect 223068 397564 223132 397628
rect 223804 397564 223868 397628
rect 225460 397564 225524 397628
rect 228772 397564 228836 397628
rect 230060 397564 230124 397628
rect 230796 397564 230860 397628
rect 232820 397564 232884 397628
rect 234292 397564 234356 397628
rect 235396 397564 235460 397628
rect 237052 397564 237116 397628
rect 238156 397564 238220 397628
rect 239628 397564 239692 397628
rect 241100 397564 241164 397628
rect 242388 397564 242452 397628
rect 243860 397564 243924 397628
rect 244596 397564 244660 397628
rect 246436 397564 246500 397628
rect 248092 397564 248156 397628
rect 248828 397564 248892 397628
rect 250852 397564 250916 397628
rect 252140 397564 252204 397628
rect 253428 397564 253492 397628
rect 254716 397564 254780 397628
rect 211292 397488 211356 397492
rect 211292 397432 211342 397488
rect 211342 397432 211356 397488
rect 211292 397428 211356 397432
rect 212580 397488 212644 397492
rect 212580 397432 212594 397488
rect 212594 397432 212644 397488
rect 212580 397428 212644 397432
rect 212764 397488 212828 397492
rect 212764 397432 212778 397488
rect 212778 397432 212828 397488
rect 212764 397428 212828 397432
rect 214236 397488 214300 397492
rect 214236 397432 214250 397488
rect 214250 397432 214300 397488
rect 214236 397428 214300 397432
rect 215340 397488 215404 397492
rect 215340 397432 215390 397488
rect 215390 397432 215404 397488
rect 215340 397428 215404 397432
rect 215708 397488 215772 397492
rect 215708 397432 215758 397488
rect 215758 397432 215772 397488
rect 215708 397428 215772 397432
rect 216812 397428 216876 397492
rect 218652 397428 218716 397492
rect 219572 397428 219636 397492
rect 221044 397488 221108 397492
rect 221044 397432 221058 397488
rect 221058 397432 221108 397488
rect 221044 397428 221108 397432
rect 222148 397428 222212 397492
rect 223988 397428 224052 397492
rect 225092 397428 225156 397492
rect 226380 397428 226444 397492
rect 228404 397428 228468 397492
rect 228956 397488 229020 397492
rect 228956 397432 228970 397488
rect 228970 397432 229020 397488
rect 228956 397428 229020 397432
rect 230244 397428 230308 397492
rect 230980 397428 231044 397492
rect 233004 397488 233068 397492
rect 233004 397432 233054 397488
rect 233054 397432 233068 397488
rect 233004 397428 233068 397432
rect 234108 397488 234172 397492
rect 234108 397432 234122 397488
rect 234122 397432 234172 397488
rect 234108 397428 234172 397432
rect 235580 397428 235644 397492
rect 237236 397428 237300 397492
rect 238340 397428 238404 397492
rect 239812 397428 239876 397492
rect 241284 397488 241348 397492
rect 241284 397432 241334 397488
rect 241334 397432 241348 397488
rect 241284 397428 241348 397432
rect 242572 397428 242636 397492
rect 244044 397488 244108 397492
rect 244044 397432 244094 397488
rect 244094 397432 244108 397488
rect 244044 397428 244108 397432
rect 245516 397488 245580 397492
rect 245516 397432 245530 397488
rect 245530 397432 245580 397488
rect 245516 397428 245580 397432
rect 246252 397428 246316 397492
rect 246804 397488 246868 397492
rect 246804 397432 246854 397488
rect 246854 397432 246868 397488
rect 246804 397428 246868 397432
rect 247908 397428 247972 397492
rect 248276 397488 248340 397492
rect 248276 397432 248290 397488
rect 248290 397432 248340 397488
rect 248276 397428 248340 397432
rect 249012 397428 249076 397492
rect 250668 397428 250732 397492
rect 252324 397488 252388 397492
rect 252324 397432 252374 397488
rect 252374 397432 252388 397488
rect 252324 397428 252388 397432
rect 253612 397488 253676 397492
rect 253612 397432 253626 397488
rect 253626 397432 253676 397488
rect 253612 397428 253676 397432
rect 254900 397428 254964 397492
rect 255268 396612 255332 396676
rect 219756 395660 219820 395724
rect 230428 395660 230492 395724
rect 215892 395524 215956 395588
rect 212580 395388 212644 395452
rect 251036 395388 251100 395452
rect 253060 395252 253124 395316
rect 226380 394300 226444 394364
rect 223068 394164 223132 394228
rect 217180 394028 217244 394092
rect 214420 393892 214484 393956
rect 235396 393892 235460 393956
rect 236868 355540 236932 355604
rect 238156 355404 238220 355468
rect 212764 355268 212828 355332
rect 248644 355268 248708 355332
rect 234108 354316 234172 354380
rect 219020 354180 219084 354244
rect 243492 354180 243556 354244
rect 215708 354044 215772 354108
rect 244596 354044 244660 354108
rect 211476 353908 211540 353972
rect 228588 353908 228652 353972
rect 253244 353908 253308 353972
rect 229876 353500 229940 353564
rect 228404 353364 228468 353428
rect 225092 352956 225156 353020
rect 237052 352956 237116 353020
rect 224172 352820 224236 352884
rect 242388 352820 242452 352884
rect 221228 352684 221292 352748
rect 247724 352684 247788 352748
rect 219572 352548 219636 352612
rect 251772 352548 251836 352612
rect 255820 351868 255884 351932
rect 222148 351324 222212 351388
rect 219940 351188 220004 351252
rect 241100 351188 241164 351252
rect 214236 351052 214300 351116
rect 251956 351052 252020 351116
rect 262628 298148 262692 298212
rect 216812 177380 216876 177444
rect 216996 177244 217060 177308
rect 232636 87620 232700 87684
rect 243676 87484 243740 87548
rect 260604 45596 260668 45660
rect 246252 26828 246316 26892
rect 237236 25468 237300 25532
rect 252140 24244 252204 24308
rect 254900 24108 254964 24172
rect 246436 22748 246500 22812
rect 248828 22612 248892 22676
rect 243860 21252 243924 21316
rect 239628 20164 239692 20228
rect 239444 20028 239508 20092
rect 246620 19892 246684 19956
rect 298508 19348 298572 19412
rect 232820 18532 232884 18596
rect 230796 17444 230860 17508
rect 253612 17308 253676 17372
rect 253428 17172 253492 17236
rect 250668 15948 250732 16012
rect 250852 15812 250916 15876
rect 246804 14724 246868 14788
rect 247908 14588 247972 14652
rect 218836 14452 218900 14516
rect 248092 14452 248156 14516
rect 216628 13228 216692 13292
rect 215524 13092 215588 13156
rect 244044 13092 244108 13156
rect 211292 12956 211356 13020
rect 245516 12956 245580 13020
rect 241284 11868 241348 11932
rect 242756 11732 242820 11796
rect 211108 11596 211172 11660
rect 242572 11596 242636 11660
rect 238340 10508 238404 10572
rect 218652 10372 218716 10436
rect 239996 10372 240060 10436
rect 215340 10236 215404 10300
rect 239812 10236 239876 10300
rect 223988 9012 224052 9076
rect 230980 9012 231044 9076
rect 214052 8876 214116 8940
rect 235580 8876 235644 8940
rect 223804 7788 223868 7852
rect 233004 7788 233068 7852
rect 220860 7652 220924 7716
rect 234292 7652 234356 7716
rect 221044 7516 221108 7580
rect 233924 7516 233988 7580
rect 224908 6156 224972 6220
rect 254716 6156 254780 6220
rect 230244 5340 230308 5404
rect 230060 5204 230124 5268
rect 237972 5068 238036 5132
rect 249012 4932 249076 4996
rect 209820 4796 209884 4860
rect 252324 4796 252388 4860
rect 226196 3708 226260 3772
rect 248276 3572 248340 3636
rect 228956 3436 229020 3500
rect 250484 3436 250548 3500
rect 223620 3300 223684 3364
rect 228772 3300 228836 3364
rect 262076 3300 262140 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 691292 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 691292 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 691292 87914 700398
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 691292 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 691292 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 691292 123914 700398
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 691292 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 691292 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 691292 159914 700398
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 80952 687454 81300 687486
rect 80952 687218 81008 687454
rect 81244 687218 81300 687454
rect 80952 687134 81300 687218
rect 80952 686898 81008 687134
rect 81244 686898 81300 687134
rect 80952 686866 81300 686898
rect 169760 687454 170108 687486
rect 169760 687218 169816 687454
rect 170052 687218 170108 687454
rect 169760 687134 170108 687218
rect 169760 686898 169816 687134
rect 170052 686898 170108 687134
rect 169760 686866 170108 686898
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 80272 655954 80620 655986
rect 80272 655718 80328 655954
rect 80564 655718 80620 655954
rect 80272 655634 80620 655718
rect 80272 655398 80328 655634
rect 80564 655398 80620 655634
rect 80272 655366 80620 655398
rect 170440 655954 170788 655986
rect 170440 655718 170496 655954
rect 170732 655718 170788 655954
rect 170440 655634 170788 655718
rect 170440 655398 170496 655634
rect 170732 655398 170788 655634
rect 170440 655366 170788 655398
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 80952 651454 81300 651486
rect 80952 651218 81008 651454
rect 81244 651218 81300 651454
rect 80952 651134 81300 651218
rect 80952 650898 81008 651134
rect 81244 650898 81300 651134
rect 80952 650866 81300 650898
rect 169760 651454 170108 651486
rect 169760 651218 169816 651454
rect 170052 651218 170108 651454
rect 169760 651134 170108 651218
rect 169760 650898 169816 651134
rect 170052 650898 170108 651134
rect 169760 650866 170108 650898
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 80272 619954 80620 619986
rect 80272 619718 80328 619954
rect 80564 619718 80620 619954
rect 80272 619634 80620 619718
rect 80272 619398 80328 619634
rect 80564 619398 80620 619634
rect 80272 619366 80620 619398
rect 170440 619954 170788 619986
rect 170440 619718 170496 619954
rect 170732 619718 170788 619954
rect 170440 619634 170788 619718
rect 170440 619398 170496 619634
rect 170732 619398 170788 619634
rect 170440 619366 170788 619398
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 80952 615454 81300 615486
rect 80952 615218 81008 615454
rect 81244 615218 81300 615454
rect 80952 615134 81300 615218
rect 80952 614898 81008 615134
rect 81244 614898 81300 615134
rect 80952 614866 81300 614898
rect 169760 615454 170108 615486
rect 169760 615218 169816 615454
rect 170052 615218 170108 615454
rect 169760 615134 170108 615218
rect 169760 614898 169816 615134
rect 170052 614898 170108 615134
rect 169760 614866 170108 614898
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 92928 599450 92988 600100
rect 94288 599450 94348 600100
rect 95376 599450 95436 600100
rect 92928 599390 93042 599450
rect 92982 597413 93042 599390
rect 94270 599390 94348 599450
rect 95374 599390 95436 599450
rect 97688 599450 97748 600100
rect 98912 599450 98972 600100
rect 100000 599450 100060 600100
rect 101088 599450 101148 600100
rect 97688 599390 97826 599450
rect 92979 597412 93045 597413
rect 92979 597348 92980 597412
rect 93044 597348 93045 597412
rect 92979 597347 93045 597348
rect 94270 597141 94330 599390
rect 94267 597140 94333 597141
rect 94267 597076 94268 597140
rect 94332 597076 94333 597140
rect 94267 597075 94333 597076
rect 95374 596325 95434 599390
rect 97766 597277 97826 599390
rect 98870 599390 98972 599450
rect 99974 599390 100060 599450
rect 101078 599390 101148 599450
rect 102312 599450 102372 600100
rect 103400 599450 103460 600100
rect 104760 599450 104820 600100
rect 102312 599390 102426 599450
rect 98870 597413 98930 599390
rect 98867 597412 98933 597413
rect 98867 597348 98868 597412
rect 98932 597348 98933 597412
rect 98867 597347 98933 597348
rect 97763 597276 97829 597277
rect 97763 597212 97764 597276
rect 97828 597212 97829 597276
rect 97763 597211 97829 597212
rect 99974 597005 100034 599390
rect 101078 597005 101138 599390
rect 102366 597549 102426 599390
rect 103286 599390 103460 599450
rect 104758 599390 104820 599450
rect 105304 599450 105364 600100
rect 105712 599450 105772 600100
rect 110472 599450 110532 600100
rect 105304 599390 105370 599450
rect 102363 597548 102429 597549
rect 102363 597484 102364 597548
rect 102428 597484 102429 597548
rect 102363 597483 102429 597484
rect 103286 597141 103346 599390
rect 103283 597140 103349 597141
rect 103283 597076 103284 597140
rect 103348 597076 103349 597140
rect 103283 597075 103349 597076
rect 99971 597004 100037 597005
rect 99971 596940 99972 597004
rect 100036 596940 100037 597004
rect 99971 596939 100037 596940
rect 101075 597004 101141 597005
rect 101075 596940 101076 597004
rect 101140 596940 101141 597004
rect 101075 596939 101141 596940
rect 104758 596869 104818 599390
rect 105310 597549 105370 599390
rect 105678 599390 105772 599450
rect 110462 599390 110532 599450
rect 115504 599450 115564 600100
rect 120536 599450 120596 600100
rect 125568 599450 125628 600100
rect 115504 599390 115674 599450
rect 120536 599390 120642 599450
rect 105307 597548 105373 597549
rect 105307 597484 105308 597548
rect 105372 597484 105373 597548
rect 105307 597483 105373 597484
rect 105678 597141 105738 599390
rect 110462 597549 110522 599390
rect 115614 597549 115674 599390
rect 120582 597549 120642 599390
rect 125550 599390 125628 599450
rect 130464 599450 130524 600100
rect 135496 599450 135556 600100
rect 130464 599390 130578 599450
rect 125550 597549 125610 599390
rect 130518 597549 130578 599390
rect 135486 599390 135556 599450
rect 140528 599450 140588 600100
rect 140528 599390 140698 599450
rect 135486 597549 135546 599390
rect 140638 597549 140698 599390
rect 106227 597548 106293 597549
rect 106227 597484 106228 597548
rect 106292 597484 106293 597548
rect 106227 597483 106293 597484
rect 110459 597548 110525 597549
rect 110459 597484 110460 597548
rect 110524 597484 110525 597548
rect 110459 597483 110525 597484
rect 115611 597548 115677 597549
rect 115611 597484 115612 597548
rect 115676 597484 115677 597548
rect 115611 597483 115677 597484
rect 120579 597548 120645 597549
rect 120579 597484 120580 597548
rect 120644 597484 120645 597548
rect 120579 597483 120645 597484
rect 125547 597548 125613 597549
rect 125547 597484 125548 597548
rect 125612 597484 125613 597548
rect 125547 597483 125613 597484
rect 130515 597548 130581 597549
rect 130515 597484 130516 597548
rect 130580 597484 130581 597548
rect 130515 597483 130581 597484
rect 135483 597548 135549 597549
rect 135483 597484 135484 597548
rect 135548 597484 135549 597548
rect 135483 597483 135549 597484
rect 140635 597548 140701 597549
rect 140635 597484 140636 597548
rect 140700 597484 140701 597548
rect 140635 597483 140701 597484
rect 105675 597140 105741 597141
rect 105675 597076 105676 597140
rect 105740 597076 105741 597140
rect 106230 597138 106290 597483
rect 106411 597140 106477 597141
rect 106411 597138 106412 597140
rect 106230 597078 106412 597138
rect 105675 597075 105741 597076
rect 106411 597076 106412 597078
rect 106476 597076 106477 597140
rect 106411 597075 106477 597076
rect 104755 596868 104821 596869
rect 104755 596804 104756 596868
rect 104820 596804 104821 596868
rect 104755 596803 104821 596804
rect 95371 596324 95437 596325
rect 95371 596260 95372 596324
rect 95436 596260 95437 596324
rect 95371 596259 95437 596260
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 80272 547954 80620 547986
rect 80272 547718 80328 547954
rect 80564 547718 80620 547954
rect 80272 547634 80620 547718
rect 80272 547398 80328 547634
rect 80564 547398 80620 547634
rect 80272 547366 80620 547398
rect 170440 547954 170788 547986
rect 170440 547718 170496 547954
rect 170732 547718 170788 547954
rect 170440 547634 170788 547718
rect 170440 547398 170496 547634
rect 170732 547398 170788 547634
rect 170440 547366 170788 547398
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 80952 543454 81300 543486
rect 80952 543218 81008 543454
rect 81244 543218 81300 543454
rect 80952 543134 81300 543218
rect 80952 542898 81008 543134
rect 81244 542898 81300 543134
rect 80952 542866 81300 542898
rect 169760 543454 170108 543486
rect 169760 543218 169816 543454
rect 170052 543218 170108 543454
rect 169760 543134 170108 543218
rect 169760 542898 169816 543134
rect 170052 542898 170108 543134
rect 169760 542866 170108 542898
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 80272 511954 80620 511986
rect 80272 511718 80328 511954
rect 80564 511718 80620 511954
rect 80272 511634 80620 511718
rect 80272 511398 80328 511634
rect 80564 511398 80620 511634
rect 80272 511366 80620 511398
rect 170440 511954 170788 511986
rect 170440 511718 170496 511954
rect 170732 511718 170788 511954
rect 170440 511634 170788 511718
rect 170440 511398 170496 511634
rect 170732 511398 170788 511634
rect 170440 511366 170788 511398
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 80952 507454 81300 507486
rect 80952 507218 81008 507454
rect 81244 507218 81300 507454
rect 80952 507134 81300 507218
rect 80952 506898 81008 507134
rect 81244 506898 81300 507134
rect 80952 506866 81300 506898
rect 169760 507454 170108 507486
rect 169760 507218 169816 507454
rect 170052 507218 170108 507454
rect 169760 507134 170108 507218
rect 169760 506898 169816 507134
rect 170052 506898 170108 507134
rect 169760 506866 170108 506898
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 92928 489930 92988 490106
rect 94288 489930 94348 490106
rect 95376 489930 95436 490106
rect 92928 489870 93042 489930
rect 92982 488477 93042 489870
rect 94270 489870 94348 489930
rect 95374 489870 95436 489930
rect 97688 489930 97748 490106
rect 98912 489930 98972 490106
rect 100000 489930 100060 490106
rect 101088 489930 101148 490106
rect 97688 489870 97826 489930
rect 94270 488477 94330 489870
rect 92979 488476 93045 488477
rect 92979 488412 92980 488476
rect 93044 488412 93045 488476
rect 92979 488411 93045 488412
rect 94267 488476 94333 488477
rect 94267 488412 94268 488476
rect 94332 488412 94333 488476
rect 94267 488411 94333 488412
rect 95374 488341 95434 489870
rect 97766 488477 97826 489870
rect 98870 489870 98972 489930
rect 99974 489870 100060 489930
rect 101078 489870 101148 489930
rect 102312 489930 102372 490106
rect 103400 489930 103460 490106
rect 104760 489930 104820 490106
rect 102312 489870 102426 489930
rect 98870 488477 98930 489870
rect 99974 488477 100034 489870
rect 101078 488477 101138 489870
rect 102366 488477 102426 489870
rect 103286 489870 103460 489930
rect 104758 489870 104820 489930
rect 105304 489930 105364 490106
rect 105712 489930 105772 490106
rect 110472 489930 110532 490106
rect 105304 489870 105370 489930
rect 97763 488476 97829 488477
rect 97763 488412 97764 488476
rect 97828 488412 97829 488476
rect 97763 488411 97829 488412
rect 98867 488476 98933 488477
rect 98867 488412 98868 488476
rect 98932 488412 98933 488476
rect 98867 488411 98933 488412
rect 99971 488476 100037 488477
rect 99971 488412 99972 488476
rect 100036 488412 100037 488476
rect 99971 488411 100037 488412
rect 101075 488476 101141 488477
rect 101075 488412 101076 488476
rect 101140 488412 101141 488476
rect 101075 488411 101141 488412
rect 102363 488476 102429 488477
rect 102363 488412 102364 488476
rect 102428 488412 102429 488476
rect 102363 488411 102429 488412
rect 95371 488340 95437 488341
rect 95371 488276 95372 488340
rect 95436 488276 95437 488340
rect 95371 488275 95437 488276
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 475954 78914 488000
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 480454 83414 488000
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 484954 87914 488000
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 453454 92414 488000
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 457954 96914 488000
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 462454 101414 488000
rect 103286 487525 103346 489870
rect 104758 488477 104818 489870
rect 105310 488477 105370 489870
rect 105678 489870 105772 489930
rect 110462 489870 110532 489930
rect 115504 489930 115564 490106
rect 120536 489930 120596 490106
rect 125568 489930 125628 490106
rect 115504 489870 115674 489930
rect 120536 489870 120642 489930
rect 105678 488477 105738 489870
rect 110462 489429 110522 489870
rect 110459 489428 110525 489429
rect 110459 489364 110460 489428
rect 110524 489364 110525 489428
rect 110459 489363 110525 489364
rect 115614 488477 115674 489870
rect 120582 488477 120642 489870
rect 125550 489870 125628 489930
rect 130464 489930 130524 490106
rect 135496 489930 135556 490106
rect 130464 489870 130578 489930
rect 125550 488477 125610 489870
rect 130518 488477 130578 489870
rect 135486 489870 135556 489930
rect 140528 489930 140588 490106
rect 140528 489870 140698 489930
rect 135486 488477 135546 489870
rect 140638 488477 140698 489870
rect 104755 488476 104821 488477
rect 104755 488412 104756 488476
rect 104820 488412 104821 488476
rect 104755 488411 104821 488412
rect 105307 488476 105373 488477
rect 105307 488412 105308 488476
rect 105372 488412 105373 488476
rect 105307 488411 105373 488412
rect 105675 488476 105741 488477
rect 105675 488412 105676 488476
rect 105740 488412 105741 488476
rect 105675 488411 105741 488412
rect 115611 488476 115677 488477
rect 115611 488412 115612 488476
rect 115676 488412 115677 488476
rect 115611 488411 115677 488412
rect 120579 488476 120645 488477
rect 120579 488412 120580 488476
rect 120644 488412 120645 488476
rect 120579 488411 120645 488412
rect 125547 488476 125613 488477
rect 125547 488412 125548 488476
rect 125612 488412 125613 488476
rect 125547 488411 125613 488412
rect 130515 488476 130581 488477
rect 130515 488412 130516 488476
rect 130580 488412 130581 488476
rect 130515 488411 130581 488412
rect 135483 488476 135549 488477
rect 135483 488412 135484 488476
rect 135548 488412 135549 488476
rect 135483 488411 135549 488412
rect 140635 488476 140701 488477
rect 140635 488412 140636 488476
rect 140700 488412 140701 488476
rect 140635 488411 140701 488412
rect 103283 487524 103349 487525
rect 103283 487460 103284 487524
rect 103348 487460 103349 487524
rect 103283 487459 103349 487460
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 466954 105914 488000
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 471454 110414 488000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 475954 114914 488000
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 480454 119414 488000
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 484954 123914 488000
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 453454 128414 488000
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 457954 132914 488000
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 462454 137414 488000
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 466954 141914 488000
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 471454 146414 488000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 475954 150914 488000
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 480454 155414 488000
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 484954 159914 488000
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 453454 164414 488000
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 457954 168914 488000
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 462454 173414 488000
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 691292 191414 695898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 691292 195914 700398
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 691292 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 691292 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 691292 231914 700398
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 691292 258914 691398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 691292 263414 695898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 691292 267914 700398
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 282131 699820 282197 699821
rect 282131 699756 282132 699820
rect 282196 699756 282197 699820
rect 282131 699755 282197 699756
rect 190952 687454 191300 687486
rect 190952 687218 191008 687454
rect 191244 687218 191300 687454
rect 190952 687134 191300 687218
rect 190952 686898 191008 687134
rect 191244 686898 191300 687134
rect 190952 686866 191300 686898
rect 279760 687454 280108 687486
rect 279760 687218 279816 687454
rect 280052 687218 280108 687454
rect 279760 687134 280108 687218
rect 279760 686898 279816 687134
rect 280052 686898 280108 687134
rect 279760 686866 280108 686898
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 190272 655954 190620 655986
rect 190272 655718 190328 655954
rect 190564 655718 190620 655954
rect 190272 655634 190620 655718
rect 190272 655398 190328 655634
rect 190564 655398 190620 655634
rect 190272 655366 190620 655398
rect 280440 655954 280788 655986
rect 280440 655718 280496 655954
rect 280732 655718 280788 655954
rect 280440 655634 280788 655718
rect 280440 655398 280496 655634
rect 280732 655398 280788 655634
rect 280440 655366 280788 655398
rect 190952 651454 191300 651486
rect 190952 651218 191008 651454
rect 191244 651218 191300 651454
rect 190952 651134 191300 651218
rect 190952 650898 191008 651134
rect 191244 650898 191300 651134
rect 190952 650866 191300 650898
rect 279760 651454 280108 651486
rect 279760 651218 279816 651454
rect 280052 651218 280108 651454
rect 279760 651134 280108 651218
rect 279760 650898 279816 651134
rect 280052 650898 280108 651134
rect 279760 650866 280108 650898
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 190272 619954 190620 619986
rect 190272 619718 190328 619954
rect 190564 619718 190620 619954
rect 190272 619634 190620 619718
rect 190272 619398 190328 619634
rect 190564 619398 190620 619634
rect 190272 619366 190620 619398
rect 280440 619954 280788 619986
rect 280440 619718 280496 619954
rect 280732 619718 280788 619954
rect 280440 619634 280788 619718
rect 280440 619398 280496 619634
rect 280732 619398 280788 619634
rect 280440 619366 280788 619398
rect 190952 615454 191300 615486
rect 190952 615218 191008 615454
rect 191244 615218 191300 615454
rect 190952 615134 191300 615218
rect 190952 614898 191008 615134
rect 191244 614898 191300 615134
rect 190952 614866 191300 614898
rect 279760 615454 280108 615486
rect 279760 615218 279816 615454
rect 280052 615218 280108 615454
rect 279760 615134 280108 615218
rect 279760 614898 279816 615134
rect 280052 614898 280108 615134
rect 279760 614866 280108 614898
rect 202928 599450 202988 600100
rect 202830 599390 202988 599450
rect 204288 599450 204348 600100
rect 205376 599450 205436 600100
rect 207688 599450 207748 600100
rect 208912 599450 208972 600100
rect 204288 599390 204362 599450
rect 205376 599390 205466 599450
rect 202830 596461 202890 599390
rect 202827 596460 202893 596461
rect 202827 596396 202828 596460
rect 202892 596396 202893 596460
rect 202827 596395 202893 596396
rect 204302 596325 204362 599390
rect 205406 596597 205466 599390
rect 207614 599390 207748 599450
rect 208902 599390 208972 599450
rect 210000 599450 210060 600100
rect 211088 599450 211148 600100
rect 212312 599450 212372 600100
rect 213400 599450 213460 600100
rect 214760 599450 214820 600100
rect 215304 599450 215364 600100
rect 215712 599450 215772 600100
rect 220472 599450 220532 600100
rect 225504 599450 225564 600100
rect 210000 599390 210066 599450
rect 211088 599390 211170 599450
rect 212312 599390 212458 599450
rect 213400 599390 213562 599450
rect 214760 599390 214850 599450
rect 215304 599390 215402 599450
rect 207614 597277 207674 599390
rect 208902 597413 208962 599390
rect 210006 597549 210066 599390
rect 210003 597548 210069 597549
rect 210003 597484 210004 597548
rect 210068 597484 210069 597548
rect 210003 597483 210069 597484
rect 208899 597412 208965 597413
rect 208899 597348 208900 597412
rect 208964 597348 208965 597412
rect 208899 597347 208965 597348
rect 207611 597276 207677 597277
rect 207611 597212 207612 597276
rect 207676 597212 207677 597276
rect 207611 597211 207677 597212
rect 211110 597005 211170 599390
rect 212398 597549 212458 599390
rect 213502 597549 213562 599390
rect 214790 597549 214850 599390
rect 212395 597548 212461 597549
rect 212395 597484 212396 597548
rect 212460 597484 212461 597548
rect 212395 597483 212461 597484
rect 213499 597548 213565 597549
rect 213499 597484 213500 597548
rect 213564 597484 213565 597548
rect 213499 597483 213565 597484
rect 214787 597548 214853 597549
rect 214787 597484 214788 597548
rect 214852 597484 214853 597548
rect 214787 597483 214853 597484
rect 215342 597141 215402 599390
rect 215710 599390 215772 599450
rect 219206 599390 220532 599450
rect 225462 599390 225564 599450
rect 230536 599450 230596 600100
rect 235568 599450 235628 600100
rect 240464 599450 240524 600100
rect 245496 599450 245556 600100
rect 250528 599450 250588 600100
rect 230536 599390 230674 599450
rect 235568 599390 235642 599450
rect 240464 599390 240610 599450
rect 245496 599390 245578 599450
rect 215710 597549 215770 599390
rect 219206 597549 219266 599390
rect 225462 597549 225522 599390
rect 230614 597549 230674 599390
rect 235582 597549 235642 599390
rect 240550 597549 240610 599390
rect 245518 597549 245578 599390
rect 250486 599390 250588 599450
rect 250486 597549 250546 599390
rect 215707 597548 215773 597549
rect 215707 597484 215708 597548
rect 215772 597484 215773 597548
rect 215707 597483 215773 597484
rect 219203 597548 219269 597549
rect 219203 597484 219204 597548
rect 219268 597484 219269 597548
rect 219203 597483 219269 597484
rect 225459 597548 225525 597549
rect 225459 597484 225460 597548
rect 225524 597484 225525 597548
rect 225459 597483 225525 597484
rect 230611 597548 230677 597549
rect 230611 597484 230612 597548
rect 230676 597484 230677 597548
rect 230611 597483 230677 597484
rect 235579 597548 235645 597549
rect 235579 597484 235580 597548
rect 235644 597484 235645 597548
rect 235579 597483 235645 597484
rect 240547 597548 240613 597549
rect 240547 597484 240548 597548
rect 240612 597484 240613 597548
rect 240547 597483 240613 597484
rect 245515 597548 245581 597549
rect 245515 597484 245516 597548
rect 245580 597484 245581 597548
rect 245515 597483 245581 597484
rect 250483 597548 250549 597549
rect 250483 597484 250484 597548
rect 250548 597484 250549 597548
rect 250483 597483 250549 597484
rect 215339 597140 215405 597141
rect 215339 597076 215340 597140
rect 215404 597076 215405 597140
rect 215339 597075 215405 597076
rect 211107 597004 211173 597005
rect 211107 596940 211108 597004
rect 211172 596940 211173 597004
rect 211107 596939 211173 596940
rect 205403 596596 205469 596597
rect 205403 596532 205404 596596
rect 205468 596532 205469 596596
rect 205403 596531 205469 596532
rect 204299 596324 204365 596325
rect 204299 596260 204300 596324
rect 204364 596260 204365 596324
rect 204299 596259 204365 596260
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 190272 547954 190620 547986
rect 190272 547718 190328 547954
rect 190564 547718 190620 547954
rect 190272 547634 190620 547718
rect 190272 547398 190328 547634
rect 190564 547398 190620 547634
rect 190272 547366 190620 547398
rect 280440 547954 280788 547986
rect 280440 547718 280496 547954
rect 280732 547718 280788 547954
rect 280440 547634 280788 547718
rect 280440 547398 280496 547634
rect 280732 547398 280788 547634
rect 280440 547366 280788 547398
rect 190952 543454 191300 543486
rect 190952 543218 191008 543454
rect 191244 543218 191300 543454
rect 190952 543134 191300 543218
rect 190952 542898 191008 543134
rect 191244 542898 191300 543134
rect 190952 542866 191300 542898
rect 279760 543454 280108 543486
rect 279760 543218 279816 543454
rect 280052 543218 280108 543454
rect 279760 543134 280108 543218
rect 279760 542898 279816 543134
rect 280052 542898 280108 543134
rect 279760 542866 280108 542898
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 190272 511954 190620 511986
rect 190272 511718 190328 511954
rect 190564 511718 190620 511954
rect 190272 511634 190620 511718
rect 190272 511398 190328 511634
rect 190564 511398 190620 511634
rect 190272 511366 190620 511398
rect 280440 511954 280788 511986
rect 280440 511718 280496 511954
rect 280732 511718 280788 511954
rect 280440 511634 280788 511718
rect 280440 511398 280496 511634
rect 280732 511398 280788 511634
rect 280440 511366 280788 511398
rect 190952 507454 191300 507486
rect 190952 507218 191008 507454
rect 191244 507218 191300 507454
rect 190952 507134 191300 507218
rect 190952 506898 191008 507134
rect 191244 506898 191300 507134
rect 190952 506866 191300 506898
rect 279760 507454 280108 507486
rect 279760 507218 279816 507454
rect 280052 507218 280108 507454
rect 279760 507134 280108 507218
rect 279760 506898 279816 507134
rect 280052 506898 280108 507134
rect 279760 506866 280108 506898
rect 202928 489930 202988 490106
rect 204288 489930 204348 490106
rect 205376 489930 205436 490106
rect 207688 489930 207748 490106
rect 208912 489930 208972 490106
rect 202928 489870 203074 489930
rect 204288 489870 204362 489930
rect 205376 489870 205466 489930
rect 203014 488069 203074 489870
rect 204302 488069 204362 489870
rect 205406 488477 205466 489870
rect 207614 489870 207748 489930
rect 208902 489870 208972 489930
rect 210000 489930 210060 490106
rect 211088 489930 211148 490106
rect 212312 489930 212372 490106
rect 213400 489930 213460 490106
rect 210000 489870 210066 489930
rect 211088 489870 211170 489930
rect 205403 488476 205469 488477
rect 205403 488412 205404 488476
rect 205468 488412 205469 488476
rect 205403 488411 205469 488412
rect 203011 488068 203077 488069
rect 203011 488004 203012 488068
rect 203076 488004 203077 488068
rect 203011 488003 203077 488004
rect 204299 488068 204365 488069
rect 204299 488004 204300 488068
rect 204364 488004 204365 488068
rect 204299 488003 204365 488004
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 480454 191414 488000
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 484954 195914 488000
rect 203014 487253 203074 488003
rect 204302 487253 204362 488003
rect 205406 487389 205466 488411
rect 205403 487388 205469 487389
rect 205403 487324 205404 487388
rect 205468 487324 205469 487388
rect 205403 487323 205469 487324
rect 207614 487253 207674 489870
rect 208902 487253 208962 489870
rect 210006 487525 210066 489870
rect 211110 487933 211170 489870
rect 212214 489870 212372 489930
rect 213318 489870 213460 489930
rect 214760 489930 214820 490106
rect 215304 489930 215364 490106
rect 215712 489930 215772 490106
rect 214760 489870 214850 489930
rect 215304 489870 215402 489930
rect 212214 488069 212274 489870
rect 212211 488068 212277 488069
rect 212211 488004 212212 488068
rect 212276 488004 212277 488068
rect 212211 488003 212277 488004
rect 211107 487932 211173 487933
rect 211107 487868 211108 487932
rect 211172 487868 211173 487932
rect 211107 487867 211173 487868
rect 213318 487525 213378 489870
rect 210003 487524 210069 487525
rect 210003 487460 210004 487524
rect 210068 487460 210069 487524
rect 210003 487459 210069 487460
rect 213315 487524 213381 487525
rect 213315 487460 213316 487524
rect 213380 487460 213381 487524
rect 213315 487459 213381 487460
rect 214790 487253 214850 489870
rect 215342 488477 215402 489870
rect 215710 489870 215772 489930
rect 220472 489930 220532 490106
rect 225504 489930 225564 490106
rect 230536 489930 230596 490106
rect 220472 489870 220554 489930
rect 215339 488476 215405 488477
rect 215339 488412 215340 488476
rect 215404 488412 215405 488476
rect 215339 488411 215405 488412
rect 215710 487253 215770 489870
rect 220494 488477 220554 489870
rect 225462 489870 225564 489930
rect 230430 489870 230596 489930
rect 235568 489930 235628 490106
rect 240464 489930 240524 490106
rect 245496 489930 245556 490106
rect 250528 489930 250588 490106
rect 235568 489870 235642 489930
rect 240464 489870 240610 489930
rect 245496 489870 245578 489930
rect 225462 488477 225522 489870
rect 230430 488477 230490 489870
rect 220491 488476 220557 488477
rect 220491 488412 220492 488476
rect 220556 488412 220557 488476
rect 220491 488411 220557 488412
rect 225459 488476 225525 488477
rect 225459 488412 225460 488476
rect 225524 488412 225525 488476
rect 225459 488411 225525 488412
rect 230427 488476 230493 488477
rect 230427 488412 230428 488476
rect 230492 488412 230493 488476
rect 230427 488411 230493 488412
rect 203011 487252 203077 487253
rect 203011 487188 203012 487252
rect 203076 487188 203077 487252
rect 203011 487187 203077 487188
rect 204299 487252 204365 487253
rect 204299 487188 204300 487252
rect 204364 487188 204365 487252
rect 204299 487187 204365 487188
rect 207611 487252 207677 487253
rect 207611 487188 207612 487252
rect 207676 487188 207677 487252
rect 207611 487187 207677 487188
rect 208899 487252 208965 487253
rect 208899 487188 208900 487252
rect 208964 487188 208965 487252
rect 208899 487187 208965 487188
rect 214787 487252 214853 487253
rect 214787 487188 214788 487252
rect 214852 487188 214853 487252
rect 214787 487187 214853 487188
rect 215707 487252 215773 487253
rect 215707 487188 215708 487252
rect 215772 487188 215773 487252
rect 215707 487187 215773 487188
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 231294 484954 231914 488000
rect 235582 487933 235642 489870
rect 240550 487933 240610 489870
rect 235579 487932 235645 487933
rect 235579 487868 235580 487932
rect 235644 487868 235645 487932
rect 235579 487867 235645 487868
rect 240547 487932 240613 487933
rect 240547 487868 240548 487932
rect 240612 487868 240613 487932
rect 240547 487867 240613 487868
rect 245518 487389 245578 489870
rect 250486 489870 250588 489930
rect 250486 487525 250546 489870
rect 250483 487524 250549 487525
rect 250483 487460 250484 487524
rect 250548 487460 250549 487524
rect 250483 487459 250549 487460
rect 245515 487388 245581 487389
rect 245515 487324 245516 487388
rect 245580 487324 245581 487388
rect 245515 487323 245581 487324
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 446000 231914 448398
rect 267294 484954 267914 488000
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 257475 446860 257541 446861
rect 257475 446796 257476 446860
rect 257540 446796 257541 446860
rect 257475 446795 257541 446796
rect 254531 446180 254597 446181
rect 254531 446116 254532 446180
rect 254596 446116 254597 446180
rect 254531 446115 254597 446116
rect 253795 444140 253861 444141
rect 253795 444076 253796 444140
rect 253860 444076 253861 444140
rect 253795 444075 253861 444076
rect 212947 443868 213013 443869
rect 212947 443804 212948 443868
rect 213012 443804 213013 443868
rect 212947 443803 213013 443804
rect 232267 443868 232333 443869
rect 232267 443804 232268 443868
rect 232332 443804 232333 443868
rect 232267 443803 232333 443804
rect 233187 443868 233253 443869
rect 233187 443804 233188 443868
rect 233252 443804 233253 443868
rect 233187 443803 233253 443804
rect 234843 443868 234909 443869
rect 234843 443804 234844 443868
rect 234908 443804 234909 443868
rect 234843 443803 234909 443804
rect 210371 443460 210437 443461
rect 210371 443396 210372 443460
rect 210436 443396 210437 443460
rect 210371 443395 210437 443396
rect 210374 443053 210434 443395
rect 210371 443052 210437 443053
rect 210371 442988 210372 443052
rect 210436 442988 210437 443052
rect 210371 442987 210437 442988
rect 212950 442237 213010 443803
rect 214235 443596 214301 443597
rect 214235 443532 214236 443596
rect 214300 443532 214301 443596
rect 214235 443531 214301 443532
rect 214238 443325 214298 443531
rect 214235 443324 214301 443325
rect 214235 443260 214236 443324
rect 214300 443260 214301 443324
rect 214235 443259 214301 443260
rect 214419 443324 214485 443325
rect 214419 443260 214420 443324
rect 214484 443260 214485 443324
rect 214419 443259 214485 443260
rect 214422 443053 214482 443259
rect 214419 443052 214485 443053
rect 214419 442988 214420 443052
rect 214484 442988 214485 443052
rect 214419 442987 214485 442988
rect 232270 442645 232330 443803
rect 232267 442644 232333 442645
rect 232267 442580 232268 442644
rect 232332 442580 232333 442644
rect 232267 442579 232333 442580
rect 233190 442509 233250 443803
rect 233187 442508 233253 442509
rect 233187 442444 233188 442508
rect 233252 442444 233253 442508
rect 233187 442443 233253 442444
rect 234846 442373 234906 443803
rect 234843 442372 234909 442373
rect 234843 442308 234844 442372
rect 234908 442308 234909 442372
rect 234843 442307 234909 442308
rect 212947 442236 213013 442237
rect 212947 442172 212948 442236
rect 213012 442172 213013 442236
rect 212947 442171 213013 442172
rect 219568 439954 219888 439986
rect 219568 439718 219610 439954
rect 219846 439718 219888 439954
rect 219568 439634 219888 439718
rect 219568 439398 219610 439634
rect 219846 439398 219888 439634
rect 219568 439366 219888 439398
rect 250288 439954 250608 439986
rect 250288 439718 250330 439954
rect 250566 439718 250608 439954
rect 250288 439634 250608 439718
rect 250288 439398 250330 439634
rect 250566 439398 250608 439634
rect 250288 439366 250608 439398
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 219568 403954 219888 403986
rect 219568 403718 219610 403954
rect 219846 403718 219888 403954
rect 219568 403634 219888 403718
rect 219568 403398 219610 403634
rect 219846 403398 219888 403634
rect 219568 403366 219888 403398
rect 250288 403954 250608 403986
rect 250288 403718 250330 403954
rect 250566 403718 250608 403954
rect 250288 403634 250608 403718
rect 250288 403398 250330 403634
rect 250566 403398 250608 403634
rect 250288 403366 250608 403398
rect 253798 399533 253858 444075
rect 253059 399532 253125 399533
rect 253059 399468 253060 399532
rect 253124 399468 253125 399532
rect 253059 399467 253125 399468
rect 253795 399532 253861 399533
rect 253795 399468 253796 399532
rect 253860 399468 253861 399532
rect 253795 399467 253861 399468
rect 217179 398852 217245 398853
rect 217179 398788 217180 398852
rect 217244 398788 217245 398852
rect 217179 398787 217245 398788
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 381454 200414 398000
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 385954 204914 398000
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 390454 209414 398000
rect 209819 397764 209885 397765
rect 209819 397700 209820 397764
rect 209884 397700 209885 397764
rect 209819 397699 209885 397700
rect 211107 397764 211173 397765
rect 211107 397700 211108 397764
rect 211172 397700 211173 397764
rect 211107 397699 211173 397700
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 209822 4861 209882 397699
rect 211110 11661 211170 397699
rect 211475 397628 211541 397629
rect 211475 397564 211476 397628
rect 211540 397564 211541 397628
rect 211475 397563 211541 397564
rect 211291 397492 211357 397493
rect 211291 397428 211292 397492
rect 211356 397428 211357 397492
rect 211291 397427 211357 397428
rect 211294 13021 211354 397427
rect 211478 353973 211538 397563
rect 212579 397492 212645 397493
rect 212579 397428 212580 397492
rect 212644 397428 212645 397492
rect 212579 397427 212645 397428
rect 212763 397492 212829 397493
rect 212763 397428 212764 397492
rect 212828 397428 212829 397492
rect 212763 397427 212829 397428
rect 212582 395453 212642 397427
rect 212579 395452 212645 395453
rect 212579 395388 212580 395452
rect 212644 395388 212645 395452
rect 212579 395387 212645 395388
rect 212766 355333 212826 397427
rect 213294 394954 213914 398000
rect 214419 397900 214485 397901
rect 214419 397836 214420 397900
rect 214484 397836 214485 397900
rect 214419 397835 214485 397836
rect 214051 397628 214117 397629
rect 214051 397564 214052 397628
rect 214116 397564 214117 397628
rect 214051 397563 214117 397564
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 212763 355332 212829 355333
rect 212763 355268 212764 355332
rect 212828 355268 212829 355332
rect 212763 355267 212829 355268
rect 211475 353972 211541 353973
rect 211475 353908 211476 353972
rect 211540 353908 211541 353972
rect 211475 353907 211541 353908
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 211291 13020 211357 13021
rect 211291 12956 211292 13020
rect 211356 12956 211357 13020
rect 211291 12955 211357 12956
rect 211107 11660 211173 11661
rect 211107 11596 211108 11660
rect 211172 11596 211173 11660
rect 211107 11595 211173 11596
rect 209819 4860 209885 4861
rect 209819 4796 209820 4860
rect 209884 4796 209885 4860
rect 209819 4795 209885 4796
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 -7066 213914 34398
rect 214054 8941 214114 397563
rect 214235 397492 214301 397493
rect 214235 397428 214236 397492
rect 214300 397428 214301 397492
rect 214235 397427 214301 397428
rect 214238 351117 214298 397427
rect 214422 393957 214482 397835
rect 215891 397764 215957 397765
rect 215891 397700 215892 397764
rect 215956 397700 215957 397764
rect 215891 397699 215957 397700
rect 216995 397764 217061 397765
rect 216995 397700 216996 397764
rect 217060 397700 217061 397764
rect 216995 397699 217061 397700
rect 215523 397628 215589 397629
rect 215523 397564 215524 397628
rect 215588 397564 215589 397628
rect 215523 397563 215589 397564
rect 215339 397492 215405 397493
rect 215339 397428 215340 397492
rect 215404 397428 215405 397492
rect 215339 397427 215405 397428
rect 214419 393956 214485 393957
rect 214419 393892 214420 393956
rect 214484 393892 214485 393956
rect 214419 393891 214485 393892
rect 214235 351116 214301 351117
rect 214235 351052 214236 351116
rect 214300 351052 214301 351116
rect 214235 351051 214301 351052
rect 215342 10301 215402 397427
rect 215526 13157 215586 397563
rect 215707 397492 215773 397493
rect 215707 397428 215708 397492
rect 215772 397428 215773 397492
rect 215707 397427 215773 397428
rect 215710 354109 215770 397427
rect 215894 395589 215954 397699
rect 216627 397628 216693 397629
rect 216627 397564 216628 397628
rect 216692 397564 216693 397628
rect 216627 397563 216693 397564
rect 215891 395588 215957 395589
rect 215891 395524 215892 395588
rect 215956 395524 215957 395588
rect 215891 395523 215957 395524
rect 215707 354108 215773 354109
rect 215707 354044 215708 354108
rect 215772 354044 215773 354108
rect 215707 354043 215773 354044
rect 216630 13293 216690 397563
rect 216811 397492 216877 397493
rect 216811 397428 216812 397492
rect 216876 397428 216877 397492
rect 216811 397427 216877 397428
rect 216814 177445 216874 397427
rect 216811 177444 216877 177445
rect 216811 177380 216812 177444
rect 216876 177380 216877 177444
rect 216811 177379 216877 177380
rect 216998 177309 217058 397699
rect 217182 394093 217242 398787
rect 226195 398036 226261 398037
rect 217179 394092 217245 394093
rect 217179 394028 217180 394092
rect 217244 394028 217245 394092
rect 217179 394027 217245 394028
rect 217794 363454 218414 398000
rect 219019 397764 219085 397765
rect 219019 397700 219020 397764
rect 219084 397700 219085 397764
rect 219019 397699 219085 397700
rect 219755 397764 219821 397765
rect 219755 397700 219756 397764
rect 219820 397700 219821 397764
rect 219755 397699 219821 397700
rect 221227 397764 221293 397765
rect 221227 397700 221228 397764
rect 221292 397700 221293 397764
rect 221227 397699 221293 397700
rect 218835 397628 218901 397629
rect 218835 397564 218836 397628
rect 218900 397564 218901 397628
rect 218835 397563 218901 397564
rect 218651 397492 218717 397493
rect 218651 397428 218652 397492
rect 218716 397428 218717 397492
rect 218651 397427 218717 397428
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 216995 177308 217061 177309
rect 216995 177244 216996 177308
rect 217060 177244 217061 177308
rect 216995 177243 217061 177244
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 216627 13292 216693 13293
rect 216627 13228 216628 13292
rect 216692 13228 216693 13292
rect 216627 13227 216693 13228
rect 215523 13156 215589 13157
rect 215523 13092 215524 13156
rect 215588 13092 215589 13156
rect 215523 13091 215589 13092
rect 215339 10300 215405 10301
rect 215339 10236 215340 10300
rect 215404 10236 215405 10300
rect 215339 10235 215405 10236
rect 214051 8940 214117 8941
rect 214051 8876 214052 8940
rect 214116 8876 214117 8940
rect 214051 8875 214117 8876
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 3454 218414 38898
rect 218654 10437 218714 397427
rect 218838 14517 218898 397563
rect 219022 354245 219082 397699
rect 219571 397492 219637 397493
rect 219571 397428 219572 397492
rect 219636 397428 219637 397492
rect 219571 397427 219637 397428
rect 219019 354244 219085 354245
rect 219019 354180 219020 354244
rect 219084 354180 219085 354244
rect 219019 354179 219085 354180
rect 219574 352613 219634 397427
rect 219758 395725 219818 397699
rect 219939 397628 220005 397629
rect 219939 397564 219940 397628
rect 220004 397564 220005 397628
rect 219939 397563 220005 397564
rect 220859 397628 220925 397629
rect 220859 397564 220860 397628
rect 220924 397564 220925 397628
rect 220859 397563 220925 397564
rect 219755 395724 219821 395725
rect 219755 395660 219756 395724
rect 219820 395660 219821 395724
rect 219755 395659 219821 395660
rect 219571 352612 219637 352613
rect 219571 352548 219572 352612
rect 219636 352548 219637 352612
rect 219571 352547 219637 352548
rect 219942 351253 220002 397563
rect 219939 351252 220005 351253
rect 219939 351188 219940 351252
rect 220004 351188 220005 351252
rect 219939 351187 220005 351188
rect 218835 14516 218901 14517
rect 218835 14452 218836 14516
rect 218900 14452 218901 14516
rect 218835 14451 218901 14452
rect 218651 10436 218717 10437
rect 218651 10372 218652 10436
rect 218716 10372 218717 10436
rect 218651 10371 218717 10372
rect 220862 7717 220922 397563
rect 221043 397492 221109 397493
rect 221043 397428 221044 397492
rect 221108 397428 221109 397492
rect 221043 397427 221109 397428
rect 220859 7716 220925 7717
rect 220859 7652 220860 7716
rect 220924 7652 220925 7716
rect 220859 7651 220925 7652
rect 221046 7581 221106 397427
rect 221230 352749 221290 397699
rect 222147 397492 222213 397493
rect 222147 397428 222148 397492
rect 222212 397428 222213 397492
rect 222147 397427 222213 397428
rect 221227 352748 221293 352749
rect 221227 352684 221228 352748
rect 221292 352684 221293 352748
rect 221227 352683 221293 352684
rect 222150 351389 222210 397427
rect 222294 367954 222914 398000
rect 226195 397972 226196 398036
rect 226260 397972 226261 398036
rect 226195 397971 226261 397972
rect 224171 397900 224237 397901
rect 224171 397836 224172 397900
rect 224236 397836 224237 397900
rect 224171 397835 224237 397836
rect 223619 397764 223685 397765
rect 223619 397700 223620 397764
rect 223684 397700 223685 397764
rect 223619 397699 223685 397700
rect 223067 397628 223133 397629
rect 223067 397564 223068 397628
rect 223132 397564 223133 397628
rect 223067 397563 223133 397564
rect 223070 394229 223130 397563
rect 223067 394228 223133 394229
rect 223067 394164 223068 394228
rect 223132 394164 223133 394228
rect 223067 394163 223133 394164
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222147 351388 222213 351389
rect 222147 351324 222148 351388
rect 222212 351324 222213 351388
rect 222147 351323 222213 351324
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 221043 7580 221109 7581
rect 221043 7516 221044 7580
rect 221108 7516 221109 7580
rect 221043 7515 221109 7516
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 223622 3365 223682 397699
rect 223803 397628 223869 397629
rect 223803 397564 223804 397628
rect 223868 397564 223869 397628
rect 223803 397563 223869 397564
rect 223806 7853 223866 397563
rect 223987 397492 224053 397493
rect 223987 397428 223988 397492
rect 224052 397428 224053 397492
rect 223987 397427 224053 397428
rect 223990 9077 224050 397427
rect 224174 352885 224234 397835
rect 225459 397628 225525 397629
rect 225459 397564 225460 397628
rect 225524 397564 225525 397628
rect 225459 397563 225525 397564
rect 225091 397492 225157 397493
rect 225091 397428 225092 397492
rect 225156 397428 225157 397492
rect 225091 397427 225157 397428
rect 225094 389330 225154 397427
rect 224910 389270 225154 389330
rect 224171 352884 224237 352885
rect 224171 352820 224172 352884
rect 224236 352820 224237 352884
rect 224171 352819 224237 352820
rect 223987 9076 224053 9077
rect 223987 9012 223988 9076
rect 224052 9012 224053 9076
rect 223987 9011 224053 9012
rect 223803 7852 223869 7853
rect 223803 7788 223804 7852
rect 223868 7788 223869 7852
rect 223803 7787 223869 7788
rect 224910 6221 224970 389270
rect 225462 389190 225522 397563
rect 225094 389130 225522 389190
rect 225094 353021 225154 389130
rect 225091 353020 225157 353021
rect 225091 352956 225092 353020
rect 225156 352956 225157 353020
rect 225091 352955 225157 352956
rect 224907 6220 224973 6221
rect 224907 6156 224908 6220
rect 224972 6156 224973 6220
rect 224907 6155 224973 6156
rect 226198 3773 226258 397971
rect 226379 397492 226445 397493
rect 226379 397428 226380 397492
rect 226444 397428 226445 397492
rect 226379 397427 226445 397428
rect 226382 394365 226442 397427
rect 226379 394364 226445 394365
rect 226379 394300 226380 394364
rect 226444 394300 226445 394364
rect 226379 394299 226445 394300
rect 226794 372454 227414 398000
rect 230427 397900 230493 397901
rect 230427 397836 230428 397900
rect 230492 397836 230493 397900
rect 230427 397835 230493 397836
rect 228587 397764 228653 397765
rect 228587 397700 228588 397764
rect 228652 397700 228653 397764
rect 228587 397699 228653 397700
rect 229875 397764 229941 397765
rect 229875 397700 229876 397764
rect 229940 397700 229941 397764
rect 229875 397699 229941 397700
rect 228403 397492 228469 397493
rect 228403 397428 228404 397492
rect 228468 397428 228469 397492
rect 228403 397427 228469 397428
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 228406 353429 228466 397427
rect 228590 353973 228650 397699
rect 228771 397628 228837 397629
rect 228771 397564 228772 397628
rect 228836 397564 228837 397628
rect 228771 397563 228837 397564
rect 228587 353972 228653 353973
rect 228587 353908 228588 353972
rect 228652 353908 228653 353972
rect 228587 353907 228653 353908
rect 228403 353428 228469 353429
rect 228403 353364 228404 353428
rect 228468 353364 228469 353428
rect 228403 353363 228469 353364
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226195 3772 226261 3773
rect 226195 3708 226196 3772
rect 226260 3708 226261 3772
rect 226195 3707 226261 3708
rect 223619 3364 223685 3365
rect 223619 3300 223620 3364
rect 223684 3300 223685 3364
rect 223619 3299 223685 3300
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 -2266 227414 11898
rect 228774 3365 228834 397563
rect 228955 397492 229021 397493
rect 228955 397428 228956 397492
rect 229020 397428 229021 397492
rect 228955 397427 229021 397428
rect 228958 3501 229018 397427
rect 229878 353565 229938 397699
rect 230059 397628 230125 397629
rect 230059 397564 230060 397628
rect 230124 397564 230125 397628
rect 230059 397563 230125 397564
rect 229875 353564 229941 353565
rect 229875 353500 229876 353564
rect 229940 353500 229941 353564
rect 229875 353499 229941 353500
rect 230062 5269 230122 397563
rect 230243 397492 230309 397493
rect 230243 397428 230244 397492
rect 230308 397428 230309 397492
rect 230243 397427 230309 397428
rect 230246 5405 230306 397427
rect 230430 395725 230490 397835
rect 230795 397628 230861 397629
rect 230795 397564 230796 397628
rect 230860 397564 230861 397628
rect 230795 397563 230861 397564
rect 230427 395724 230493 395725
rect 230427 395660 230428 395724
rect 230492 395660 230493 395724
rect 230427 395659 230493 395660
rect 230798 17509 230858 397563
rect 230979 397492 231045 397493
rect 230979 397428 230980 397492
rect 231044 397428 231045 397492
rect 230979 397427 231045 397428
rect 230795 17508 230861 17509
rect 230795 17444 230796 17508
rect 230860 17444 230861 17508
rect 230795 17443 230861 17444
rect 230982 9077 231042 397427
rect 231294 376954 231914 398000
rect 232635 397764 232701 397765
rect 232635 397700 232636 397764
rect 232700 397700 232701 397764
rect 232635 397699 232701 397700
rect 233923 397764 233989 397765
rect 233923 397700 233924 397764
rect 233988 397700 233989 397764
rect 233923 397699 233989 397700
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 232638 87685 232698 397699
rect 232819 397628 232885 397629
rect 232819 397564 232820 397628
rect 232884 397564 232885 397628
rect 232819 397563 232885 397564
rect 232635 87684 232701 87685
rect 232635 87620 232636 87684
rect 232700 87620 232701 87684
rect 232635 87619 232701 87620
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 232822 18597 232882 397563
rect 233003 397492 233069 397493
rect 233003 397428 233004 397492
rect 233068 397428 233069 397492
rect 233003 397427 233069 397428
rect 232819 18596 232885 18597
rect 232819 18532 232820 18596
rect 232884 18532 232885 18596
rect 232819 18531 232885 18532
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 230979 9076 231045 9077
rect 230979 9012 230980 9076
rect 231044 9012 231045 9076
rect 230979 9011 231045 9012
rect 230243 5404 230309 5405
rect 230243 5340 230244 5404
rect 230308 5340 230309 5404
rect 230243 5339 230309 5340
rect 230059 5268 230125 5269
rect 230059 5204 230060 5268
rect 230124 5204 230125 5268
rect 230059 5203 230125 5204
rect 228955 3500 229021 3501
rect 228955 3436 228956 3500
rect 229020 3436 229021 3500
rect 228955 3435 229021 3436
rect 228771 3364 228837 3365
rect 228771 3300 228772 3364
rect 228836 3300 228837 3364
rect 228771 3299 228837 3300
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 -3226 231914 16398
rect 233006 7853 233066 397427
rect 233003 7852 233069 7853
rect 233003 7788 233004 7852
rect 233068 7788 233069 7852
rect 233003 7787 233069 7788
rect 233926 7581 233986 397699
rect 234291 397628 234357 397629
rect 234291 397564 234292 397628
rect 234356 397564 234357 397628
rect 234291 397563 234357 397564
rect 235395 397628 235461 397629
rect 235395 397564 235396 397628
rect 235460 397564 235461 397628
rect 235395 397563 235461 397564
rect 234107 397492 234173 397493
rect 234107 397428 234108 397492
rect 234172 397428 234173 397492
rect 234107 397427 234173 397428
rect 234110 354381 234170 397427
rect 234107 354380 234173 354381
rect 234107 354316 234108 354380
rect 234172 354316 234173 354380
rect 234107 354315 234173 354316
rect 234294 7717 234354 397563
rect 235398 393957 235458 397563
rect 235579 397492 235645 397493
rect 235579 397428 235580 397492
rect 235644 397428 235645 397492
rect 235579 397427 235645 397428
rect 235395 393956 235461 393957
rect 235395 393892 235396 393956
rect 235460 393892 235461 393956
rect 235395 393891 235461 393892
rect 235582 8941 235642 397427
rect 235794 381454 236414 398000
rect 239443 397900 239509 397901
rect 239443 397836 239444 397900
rect 239508 397836 239509 397900
rect 239443 397835 239509 397836
rect 236867 397764 236933 397765
rect 236867 397700 236868 397764
rect 236932 397700 236933 397764
rect 236867 397699 236933 397700
rect 237971 397764 238037 397765
rect 237971 397700 237972 397764
rect 238036 397700 238037 397764
rect 237971 397699 238037 397700
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 236870 355605 236930 397699
rect 237051 397628 237117 397629
rect 237051 397564 237052 397628
rect 237116 397564 237117 397628
rect 237051 397563 237117 397564
rect 236867 355604 236933 355605
rect 236867 355540 236868 355604
rect 236932 355540 236933 355604
rect 236867 355539 236933 355540
rect 237054 353021 237114 397563
rect 237235 397492 237301 397493
rect 237235 397428 237236 397492
rect 237300 397428 237301 397492
rect 237235 397427 237301 397428
rect 237051 353020 237117 353021
rect 237051 352956 237052 353020
rect 237116 352956 237117 353020
rect 237051 352955 237117 352956
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 237238 25533 237298 397427
rect 237235 25532 237301 25533
rect 237235 25468 237236 25532
rect 237300 25468 237301 25532
rect 237235 25467 237301 25468
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235579 8940 235645 8941
rect 235579 8876 235580 8940
rect 235644 8876 235645 8940
rect 235579 8875 235645 8876
rect 234291 7716 234357 7717
rect 234291 7652 234292 7716
rect 234356 7652 234357 7716
rect 234291 7651 234357 7652
rect 233923 7580 233989 7581
rect 233923 7516 233924 7580
rect 233988 7516 233989 7580
rect 233923 7515 233989 7516
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 -4186 236414 20898
rect 237974 5133 238034 397699
rect 238155 397628 238221 397629
rect 238155 397564 238156 397628
rect 238220 397564 238221 397628
rect 238155 397563 238221 397564
rect 238158 355469 238218 397563
rect 238339 397492 238405 397493
rect 238339 397428 238340 397492
rect 238404 397428 238405 397492
rect 238339 397427 238405 397428
rect 238155 355468 238221 355469
rect 238155 355404 238156 355468
rect 238220 355404 238221 355468
rect 238155 355403 238221 355404
rect 238342 10573 238402 397427
rect 239446 20093 239506 397835
rect 239995 397764 240061 397765
rect 239995 397700 239996 397764
rect 240060 397700 240061 397764
rect 239995 397699 240061 397700
rect 239627 397628 239693 397629
rect 239627 397564 239628 397628
rect 239692 397564 239693 397628
rect 239627 397563 239693 397564
rect 239630 20229 239690 397563
rect 239811 397492 239877 397493
rect 239811 397428 239812 397492
rect 239876 397428 239877 397492
rect 239811 397427 239877 397428
rect 239627 20228 239693 20229
rect 239627 20164 239628 20228
rect 239692 20164 239693 20228
rect 239627 20163 239693 20164
rect 239443 20092 239509 20093
rect 239443 20028 239444 20092
rect 239508 20028 239509 20092
rect 239443 20027 239509 20028
rect 238339 10572 238405 10573
rect 238339 10508 238340 10572
rect 238404 10508 238405 10572
rect 238339 10507 238405 10508
rect 239814 10301 239874 397427
rect 239998 10437 240058 397699
rect 240294 385954 240914 398000
rect 243491 397900 243557 397901
rect 243491 397836 243492 397900
rect 243556 397836 243557 397900
rect 243491 397835 243557 397836
rect 242755 397764 242821 397765
rect 242755 397700 242756 397764
rect 242820 397700 242821 397764
rect 242755 397699 242821 397700
rect 241099 397628 241165 397629
rect 241099 397564 241100 397628
rect 241164 397564 241165 397628
rect 241099 397563 241165 397564
rect 242387 397628 242453 397629
rect 242387 397564 242388 397628
rect 242452 397564 242453 397628
rect 242387 397563 242453 397564
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 241102 351253 241162 397563
rect 241283 397492 241349 397493
rect 241283 397428 241284 397492
rect 241348 397428 241349 397492
rect 241283 397427 241349 397428
rect 241099 351252 241165 351253
rect 241099 351188 241100 351252
rect 241164 351188 241165 351252
rect 241099 351187 241165 351188
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 239995 10436 240061 10437
rect 239995 10372 239996 10436
rect 240060 10372 240061 10436
rect 239995 10371 240061 10372
rect 239811 10300 239877 10301
rect 239811 10236 239812 10300
rect 239876 10236 239877 10300
rect 239811 10235 239877 10236
rect 237971 5132 238037 5133
rect 237971 5068 237972 5132
rect 238036 5068 238037 5132
rect 237971 5067 238037 5068
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 -5146 240914 25398
rect 241286 11933 241346 397427
rect 242390 352885 242450 397563
rect 242571 397492 242637 397493
rect 242571 397428 242572 397492
rect 242636 397428 242637 397492
rect 242571 397427 242637 397428
rect 242387 352884 242453 352885
rect 242387 352820 242388 352884
rect 242452 352820 242453 352884
rect 242387 352819 242453 352820
rect 241283 11932 241349 11933
rect 241283 11868 241284 11932
rect 241348 11868 241349 11932
rect 241283 11867 241349 11868
rect 242574 11661 242634 397427
rect 242758 11797 242818 397699
rect 243494 354245 243554 397835
rect 243675 397764 243741 397765
rect 243675 397700 243676 397764
rect 243740 397700 243741 397764
rect 243675 397699 243741 397700
rect 243491 354244 243557 354245
rect 243491 354180 243492 354244
rect 243556 354180 243557 354244
rect 243491 354179 243557 354180
rect 243678 87549 243738 397699
rect 243859 397628 243925 397629
rect 243859 397564 243860 397628
rect 243924 397564 243925 397628
rect 243859 397563 243925 397564
rect 244595 397628 244661 397629
rect 244595 397564 244596 397628
rect 244660 397564 244661 397628
rect 244595 397563 244661 397564
rect 243675 87548 243741 87549
rect 243675 87484 243676 87548
rect 243740 87484 243741 87548
rect 243675 87483 243741 87484
rect 243862 21317 243922 397563
rect 244043 397492 244109 397493
rect 244043 397428 244044 397492
rect 244108 397428 244109 397492
rect 244043 397427 244109 397428
rect 243859 21316 243925 21317
rect 243859 21252 243860 21316
rect 243924 21252 243925 21316
rect 243859 21251 243925 21252
rect 244046 13157 244106 397427
rect 244598 354109 244658 397563
rect 244794 390454 245414 398000
rect 246619 397764 246685 397765
rect 246619 397700 246620 397764
rect 246684 397700 246685 397764
rect 246619 397699 246685 397700
rect 247723 397764 247789 397765
rect 247723 397700 247724 397764
rect 247788 397700 247789 397764
rect 247723 397699 247789 397700
rect 248643 397764 248709 397765
rect 248643 397700 248644 397764
rect 248708 397700 248709 397764
rect 248643 397699 248709 397700
rect 246435 397628 246501 397629
rect 246435 397564 246436 397628
rect 246500 397564 246501 397628
rect 246435 397563 246501 397564
rect 245515 397492 245581 397493
rect 245515 397428 245516 397492
rect 245580 397428 245581 397492
rect 245515 397427 245581 397428
rect 246251 397492 246317 397493
rect 246251 397428 246252 397492
rect 246316 397428 246317 397492
rect 246251 397427 246317 397428
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244595 354108 244661 354109
rect 244595 354044 244596 354108
rect 244660 354044 244661 354108
rect 244595 354043 244661 354044
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244043 13156 244109 13157
rect 244043 13092 244044 13156
rect 244108 13092 244109 13156
rect 244043 13091 244109 13092
rect 242755 11796 242821 11797
rect 242755 11732 242756 11796
rect 242820 11732 242821 11796
rect 242755 11731 242821 11732
rect 242571 11660 242637 11661
rect 242571 11596 242572 11660
rect 242636 11596 242637 11660
rect 242571 11595 242637 11596
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 -6106 245414 29898
rect 245518 13021 245578 397427
rect 246254 26893 246314 397427
rect 246251 26892 246317 26893
rect 246251 26828 246252 26892
rect 246316 26828 246317 26892
rect 246251 26827 246317 26828
rect 246438 22813 246498 397563
rect 246435 22812 246501 22813
rect 246435 22748 246436 22812
rect 246500 22748 246501 22812
rect 246435 22747 246501 22748
rect 246622 19957 246682 397699
rect 246803 397492 246869 397493
rect 246803 397428 246804 397492
rect 246868 397428 246869 397492
rect 246803 397427 246869 397428
rect 246619 19956 246685 19957
rect 246619 19892 246620 19956
rect 246684 19892 246685 19956
rect 246619 19891 246685 19892
rect 246806 14789 246866 397427
rect 247726 352749 247786 397699
rect 248091 397628 248157 397629
rect 248091 397564 248092 397628
rect 248156 397564 248157 397628
rect 248091 397563 248157 397564
rect 247907 397492 247973 397493
rect 247907 397428 247908 397492
rect 247972 397428 247973 397492
rect 247907 397427 247973 397428
rect 247723 352748 247789 352749
rect 247723 352684 247724 352748
rect 247788 352684 247789 352748
rect 247723 352683 247789 352684
rect 246803 14788 246869 14789
rect 246803 14724 246804 14788
rect 246868 14724 246869 14788
rect 246803 14723 246869 14724
rect 247910 14653 247970 397427
rect 247907 14652 247973 14653
rect 247907 14588 247908 14652
rect 247972 14588 247973 14652
rect 247907 14587 247973 14588
rect 248094 14517 248154 397563
rect 248275 397492 248341 397493
rect 248275 397428 248276 397492
rect 248340 397428 248341 397492
rect 248275 397427 248341 397428
rect 248091 14516 248157 14517
rect 248091 14452 248092 14516
rect 248156 14452 248157 14516
rect 248091 14451 248157 14452
rect 245515 13020 245581 13021
rect 245515 12956 245516 13020
rect 245580 12956 245581 13020
rect 245515 12955 245581 12956
rect 248278 3637 248338 397427
rect 248646 355333 248706 397699
rect 248827 397628 248893 397629
rect 248827 397564 248828 397628
rect 248892 397564 248893 397628
rect 248827 397563 248893 397564
rect 248643 355332 248709 355333
rect 248643 355268 248644 355332
rect 248708 355268 248709 355332
rect 248643 355267 248709 355268
rect 248830 22677 248890 397563
rect 249011 397492 249077 397493
rect 249011 397428 249012 397492
rect 249076 397428 249077 397492
rect 249011 397427 249077 397428
rect 248827 22676 248893 22677
rect 248827 22612 248828 22676
rect 248892 22612 248893 22676
rect 248827 22611 248893 22612
rect 249014 4997 249074 397427
rect 249294 394954 249914 398000
rect 251035 397900 251101 397901
rect 251035 397836 251036 397900
rect 251100 397836 251101 397900
rect 251035 397835 251101 397836
rect 251771 397900 251837 397901
rect 251771 397836 251772 397900
rect 251836 397836 251837 397900
rect 251771 397835 251837 397836
rect 250483 397764 250549 397765
rect 250483 397700 250484 397764
rect 250548 397700 250549 397764
rect 250483 397699 250549 397700
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249011 4996 249077 4997
rect 249011 4932 249012 4996
rect 249076 4932 249077 4996
rect 249011 4931 249077 4932
rect 248275 3636 248341 3637
rect 248275 3572 248276 3636
rect 248340 3572 248341 3636
rect 248275 3571 248341 3572
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 -7066 249914 34398
rect 250486 3501 250546 397699
rect 250851 397628 250917 397629
rect 250851 397564 250852 397628
rect 250916 397564 250917 397628
rect 250851 397563 250917 397564
rect 250667 397492 250733 397493
rect 250667 397428 250668 397492
rect 250732 397428 250733 397492
rect 250667 397427 250733 397428
rect 250670 16013 250730 397427
rect 250667 16012 250733 16013
rect 250667 15948 250668 16012
rect 250732 15948 250733 16012
rect 250667 15947 250733 15948
rect 250854 15877 250914 397563
rect 251038 395453 251098 397835
rect 251035 395452 251101 395453
rect 251035 395388 251036 395452
rect 251100 395388 251101 395452
rect 251035 395387 251101 395388
rect 251774 352613 251834 397835
rect 251955 397764 252021 397765
rect 251955 397700 251956 397764
rect 252020 397700 252021 397764
rect 251955 397699 252021 397700
rect 251771 352612 251837 352613
rect 251771 352548 251772 352612
rect 251836 352548 251837 352612
rect 251771 352547 251837 352548
rect 251958 351117 252018 397699
rect 252139 397628 252205 397629
rect 252139 397564 252140 397628
rect 252204 397564 252205 397628
rect 252139 397563 252205 397564
rect 251955 351116 252021 351117
rect 251955 351052 251956 351116
rect 252020 351052 252021 351116
rect 251955 351051 252021 351052
rect 252142 24309 252202 397563
rect 252323 397492 252389 397493
rect 252323 397428 252324 397492
rect 252388 397428 252389 397492
rect 252323 397427 252389 397428
rect 252139 24308 252205 24309
rect 252139 24244 252140 24308
rect 252204 24244 252205 24308
rect 252139 24243 252205 24244
rect 250851 15876 250917 15877
rect 250851 15812 250852 15876
rect 250916 15812 250917 15876
rect 250851 15811 250917 15812
rect 252326 4861 252386 397427
rect 253062 395317 253122 399467
rect 253243 399396 253309 399397
rect 253243 399332 253244 399396
rect 253308 399332 253309 399396
rect 253243 399331 253309 399332
rect 253246 398717 253306 399331
rect 254534 399125 254594 446115
rect 257291 445772 257357 445773
rect 257291 445708 257292 445772
rect 257356 445708 257357 445772
rect 257291 445707 257357 445708
rect 254899 445636 254965 445637
rect 254899 445572 254900 445636
rect 254964 445572 254965 445636
rect 254899 445571 254965 445572
rect 254715 445092 254781 445093
rect 254715 445028 254716 445092
rect 254780 445028 254781 445092
rect 254715 445027 254781 445028
rect 254531 399124 254597 399125
rect 254531 399060 254532 399124
rect 254596 399060 254597 399124
rect 254531 399059 254597 399060
rect 253243 398716 253309 398717
rect 253243 398652 253244 398716
rect 253308 398652 253309 398716
rect 253243 398651 253309 398652
rect 253243 397764 253309 397765
rect 253243 397700 253244 397764
rect 253308 397700 253309 397764
rect 253243 397699 253309 397700
rect 253059 395316 253125 395317
rect 253059 395252 253060 395316
rect 253124 395252 253125 395316
rect 253059 395251 253125 395252
rect 253246 353973 253306 397699
rect 253427 397628 253493 397629
rect 253427 397564 253428 397628
rect 253492 397564 253493 397628
rect 253427 397563 253493 397564
rect 253243 353972 253309 353973
rect 253243 353908 253244 353972
rect 253308 353908 253309 353972
rect 253243 353907 253309 353908
rect 253430 17237 253490 397563
rect 253611 397492 253677 397493
rect 253611 397428 253612 397492
rect 253676 397428 253677 397492
rect 253611 397427 253677 397428
rect 253614 17373 253674 397427
rect 253794 363454 254414 398000
rect 254718 397901 254778 445027
rect 254902 398989 254962 445571
rect 255819 443596 255885 443597
rect 255819 443532 255820 443596
rect 255884 443532 255885 443596
rect 255819 443531 255885 443532
rect 256555 443596 256621 443597
rect 256555 443532 256556 443596
rect 256620 443532 256621 443596
rect 256555 443531 256621 443532
rect 255267 399260 255333 399261
rect 255267 399196 255268 399260
rect 255332 399196 255333 399260
rect 255267 399195 255333 399196
rect 254899 398988 254965 398989
rect 254899 398924 254900 398988
rect 254964 398924 254965 398988
rect 254899 398923 254965 398924
rect 254715 397900 254781 397901
rect 254715 397836 254716 397900
rect 254780 397836 254781 397900
rect 254715 397835 254781 397836
rect 254715 397628 254781 397629
rect 254715 397564 254716 397628
rect 254780 397564 254781 397628
rect 254715 397563 254781 397564
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253611 17372 253677 17373
rect 253611 17308 253612 17372
rect 253676 17308 253677 17372
rect 253611 17307 253677 17308
rect 253427 17236 253493 17237
rect 253427 17172 253428 17236
rect 253492 17172 253493 17236
rect 253427 17171 253493 17172
rect 252323 4860 252389 4861
rect 252323 4796 252324 4860
rect 252388 4796 252389 4860
rect 252323 4795 252389 4796
rect 250483 3500 250549 3501
rect 250483 3436 250484 3500
rect 250548 3436 250549 3500
rect 250483 3435 250549 3436
rect 253794 3454 254414 38898
rect 254718 6221 254778 397563
rect 254899 397492 254965 397493
rect 254899 397428 254900 397492
rect 254964 397428 254965 397492
rect 254899 397427 254965 397428
rect 254902 24173 254962 397427
rect 255270 396677 255330 399195
rect 255267 396676 255333 396677
rect 255267 396612 255268 396676
rect 255332 396612 255333 396676
rect 255267 396611 255333 396612
rect 255822 351933 255882 443531
rect 256558 400213 256618 443531
rect 256555 400212 256621 400213
rect 256555 400148 256556 400212
rect 256620 400148 256621 400212
rect 256555 400147 256621 400148
rect 257294 398445 257354 445707
rect 257478 399125 257538 446795
rect 262627 446724 262693 446725
rect 262627 446660 262628 446724
rect 262692 446660 262693 446724
rect 262627 446659 262693 446660
rect 260603 445636 260669 445637
rect 260603 445572 260604 445636
rect 260668 445572 260669 445636
rect 260603 445571 260669 445572
rect 260051 444412 260117 444413
rect 260051 444348 260052 444412
rect 260116 444348 260117 444412
rect 260051 444347 260117 444348
rect 259131 443460 259197 443461
rect 259131 443396 259132 443460
rect 259196 443396 259197 443460
rect 259131 443395 259197 443396
rect 259315 443460 259381 443461
rect 259315 443396 259316 443460
rect 259380 443396 259381 443460
rect 259315 443395 259381 443396
rect 259134 401573 259194 443395
rect 259131 401572 259197 401573
rect 259131 401508 259132 401572
rect 259196 401508 259197 401572
rect 259131 401507 259197 401508
rect 257475 399124 257541 399125
rect 257475 399060 257476 399124
rect 257540 399060 257541 399124
rect 257475 399059 257541 399060
rect 257291 398444 257357 398445
rect 257291 398380 257292 398444
rect 257356 398380 257357 398444
rect 257291 398379 257357 398380
rect 259318 398309 259378 443395
rect 260054 398581 260114 444347
rect 260051 398580 260117 398581
rect 260051 398516 260052 398580
rect 260116 398516 260117 398580
rect 260051 398515 260117 398516
rect 259315 398308 259381 398309
rect 259315 398244 259316 398308
rect 259380 398244 259381 398308
rect 259315 398243 259381 398244
rect 258294 367954 258914 398000
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 255819 351932 255885 351933
rect 255819 351868 255820 351932
rect 255884 351868 255885 351932
rect 255819 351867 255885 351868
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 260606 45661 260666 445571
rect 262075 443460 262141 443461
rect 262075 443396 262076 443460
rect 262140 443396 262141 443460
rect 262075 443395 262141 443396
rect 260603 45660 260669 45661
rect 260603 45596 260604 45660
rect 260668 45596 260669 45660
rect 260603 45595 260669 45596
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 254899 24172 254965 24173
rect 254899 24108 254900 24172
rect 254964 24108 254965 24172
rect 254899 24107 254965 24108
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 254715 6220 254781 6221
rect 254715 6156 254716 6220
rect 254780 6156 254781 6220
rect 254715 6155 254781 6156
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 -1306 258914 7398
rect 262078 3365 262138 443395
rect 262630 298213 262690 446659
rect 267294 446000 267914 448398
rect 271794 453454 272414 488000
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 263547 398444 263613 398445
rect 263547 398380 263548 398444
rect 263612 398380 263613 398444
rect 263547 398379 263613 398380
rect 262794 372454 263414 398000
rect 263550 397901 263610 398379
rect 263547 397900 263613 397901
rect 263547 397836 263548 397900
rect 263612 397836 263613 397900
rect 263547 397835 263613 397836
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262627 298212 262693 298213
rect 262627 298148 262628 298212
rect 262692 298148 262693 298212
rect 262627 298147 262693 298148
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262075 3364 262141 3365
rect 262075 3300 262076 3364
rect 262140 3300 262141 3364
rect 262075 3299 262141 3300
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 376954 267914 398000
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 457954 276914 488000
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 462454 281414 488000
rect 282134 476781 282194 699755
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 282131 476780 282197 476781
rect 282131 476716 282132 476780
rect 282196 476716 282197 476780
rect 282131 476715 282197 476716
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 691292 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 691292 303914 700398
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 691292 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 691292 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 691292 339914 700398
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 691292 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 691292 371414 695898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 691292 375914 700398
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 300952 687454 301300 687486
rect 300952 687218 301008 687454
rect 301244 687218 301300 687454
rect 300952 687134 301300 687218
rect 300952 686898 301008 687134
rect 301244 686898 301300 687134
rect 300952 686866 301300 686898
rect 389760 687454 390108 687486
rect 389760 687218 389816 687454
rect 390052 687218 390108 687454
rect 389760 687134 390108 687218
rect 389760 686898 389816 687134
rect 390052 686898 390108 687134
rect 389760 686866 390108 686898
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 300272 655954 300620 655986
rect 300272 655718 300328 655954
rect 300564 655718 300620 655954
rect 300272 655634 300620 655718
rect 300272 655398 300328 655634
rect 300564 655398 300620 655634
rect 300272 655366 300620 655398
rect 390440 655954 390788 655986
rect 390440 655718 390496 655954
rect 390732 655718 390788 655954
rect 390440 655634 390788 655718
rect 390440 655398 390496 655634
rect 390732 655398 390788 655634
rect 390440 655366 390788 655398
rect 300952 651454 301300 651486
rect 300952 651218 301008 651454
rect 301244 651218 301300 651454
rect 300952 651134 301300 651218
rect 300952 650898 301008 651134
rect 301244 650898 301300 651134
rect 300952 650866 301300 650898
rect 389760 651454 390108 651486
rect 389760 651218 389816 651454
rect 390052 651218 390108 651454
rect 389760 651134 390108 651218
rect 389760 650898 389816 651134
rect 390052 650898 390108 651134
rect 389760 650866 390108 650898
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 300272 619954 300620 619986
rect 300272 619718 300328 619954
rect 300564 619718 300620 619954
rect 300272 619634 300620 619718
rect 300272 619398 300328 619634
rect 300564 619398 300620 619634
rect 300272 619366 300620 619398
rect 390440 619954 390788 619986
rect 390440 619718 390496 619954
rect 390732 619718 390788 619954
rect 390440 619634 390788 619718
rect 390440 619398 390496 619634
rect 390732 619398 390788 619634
rect 390440 619366 390788 619398
rect 300952 615454 301300 615486
rect 300952 615218 301008 615454
rect 301244 615218 301300 615454
rect 300952 615134 301300 615218
rect 300952 614898 301008 615134
rect 301244 614898 301300 615134
rect 300952 614866 301300 614898
rect 389760 615454 390108 615486
rect 389760 615218 389816 615454
rect 390052 615218 390108 615454
rect 389760 615134 390108 615218
rect 389760 614898 389816 615134
rect 390052 614898 390108 615134
rect 389760 614866 390108 614898
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 312928 599450 312988 600100
rect 312862 599390 312988 599450
rect 314288 599450 314348 600100
rect 315376 599450 315436 600100
rect 317688 599450 317748 600100
rect 314288 599390 314394 599450
rect 312862 596325 312922 599390
rect 314334 596325 314394 599390
rect 315254 599390 315436 599450
rect 317646 599390 317748 599450
rect 318912 599450 318972 600100
rect 320000 599450 320060 600100
rect 321088 599450 321148 600100
rect 322312 599450 322372 600100
rect 323400 599450 323460 600100
rect 318912 599390 318994 599450
rect 320000 599390 320098 599450
rect 321088 599390 321202 599450
rect 315254 597413 315314 599390
rect 315251 597412 315317 597413
rect 315251 597348 315252 597412
rect 315316 597348 315317 597412
rect 315251 597347 315317 597348
rect 317646 597141 317706 599390
rect 318934 597277 318994 599390
rect 320038 597549 320098 599390
rect 320035 597548 320101 597549
rect 320035 597484 320036 597548
rect 320100 597484 320101 597548
rect 320035 597483 320101 597484
rect 321142 597413 321202 599390
rect 322246 599390 322372 599450
rect 323350 599390 323460 599450
rect 324760 599450 324820 600100
rect 325304 599450 325364 600100
rect 325712 599450 325772 600100
rect 330472 599450 330532 600100
rect 335504 599450 335564 600100
rect 340536 599450 340596 600100
rect 324760 599390 324882 599450
rect 325304 599390 325434 599450
rect 325712 599390 325802 599450
rect 330472 599390 330586 599450
rect 322246 597549 322306 599390
rect 323350 597549 323410 599390
rect 324822 597549 324882 599390
rect 322243 597548 322309 597549
rect 322243 597484 322244 597548
rect 322308 597484 322309 597548
rect 322243 597483 322309 597484
rect 323347 597548 323413 597549
rect 323347 597484 323348 597548
rect 323412 597484 323413 597548
rect 323347 597483 323413 597484
rect 324819 597548 324885 597549
rect 324819 597484 324820 597548
rect 324884 597484 324885 597548
rect 324819 597483 324885 597484
rect 321139 597412 321205 597413
rect 321139 597348 321140 597412
rect 321204 597348 321205 597412
rect 321139 597347 321205 597348
rect 318931 597276 318997 597277
rect 318931 597212 318932 597276
rect 318996 597212 318997 597276
rect 318931 597211 318997 597212
rect 317643 597140 317709 597141
rect 317643 597076 317644 597140
rect 317708 597076 317709 597140
rect 317643 597075 317709 597076
rect 321142 597005 321202 597347
rect 321139 597004 321205 597005
rect 321139 596940 321140 597004
rect 321204 596940 321205 597004
rect 321139 596939 321205 596940
rect 325374 596869 325434 599390
rect 325742 597549 325802 599390
rect 330526 597549 330586 599390
rect 335126 599390 335564 599450
rect 340462 599390 340596 599450
rect 345568 599450 345628 600100
rect 350464 599450 350524 600100
rect 355496 599450 355556 600100
rect 360528 599450 360588 600100
rect 345568 599390 345674 599450
rect 335126 597549 335186 599390
rect 340462 597549 340522 599390
rect 345614 597549 345674 599390
rect 350398 599390 350524 599450
rect 354446 599390 355556 599450
rect 360518 599390 360588 599450
rect 350398 597549 350458 599390
rect 354446 597549 354506 599390
rect 360518 597549 360578 599390
rect 325739 597548 325805 597549
rect 325739 597484 325740 597548
rect 325804 597484 325805 597548
rect 325739 597483 325805 597484
rect 330523 597548 330589 597549
rect 330523 597484 330524 597548
rect 330588 597484 330589 597548
rect 330523 597483 330589 597484
rect 335123 597548 335189 597549
rect 335123 597484 335124 597548
rect 335188 597484 335189 597548
rect 335123 597483 335189 597484
rect 340459 597548 340525 597549
rect 340459 597484 340460 597548
rect 340524 597484 340525 597548
rect 340459 597483 340525 597484
rect 345611 597548 345677 597549
rect 345611 597484 345612 597548
rect 345676 597484 345677 597548
rect 345611 597483 345677 597484
rect 350395 597548 350461 597549
rect 350395 597484 350396 597548
rect 350460 597484 350461 597548
rect 350395 597483 350461 597484
rect 354443 597548 354509 597549
rect 354443 597484 354444 597548
rect 354508 597484 354509 597548
rect 354443 597483 354509 597484
rect 360515 597548 360581 597549
rect 360515 597484 360516 597548
rect 360580 597484 360581 597548
rect 360515 597483 360581 597484
rect 325371 596868 325437 596869
rect 325371 596804 325372 596868
rect 325436 596804 325437 596868
rect 325371 596803 325437 596804
rect 312859 596324 312925 596325
rect 312859 596260 312860 596324
rect 312924 596260 312925 596324
rect 312859 596259 312925 596260
rect 314331 596324 314397 596325
rect 314331 596260 314332 596324
rect 314396 596260 314397 596324
rect 314331 596259 314397 596260
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 300272 547954 300620 547986
rect 300272 547718 300328 547954
rect 300564 547718 300620 547954
rect 300272 547634 300620 547718
rect 300272 547398 300328 547634
rect 300564 547398 300620 547634
rect 300272 547366 300620 547398
rect 390440 547954 390788 547986
rect 390440 547718 390496 547954
rect 390732 547718 390788 547954
rect 390440 547634 390788 547718
rect 390440 547398 390496 547634
rect 390732 547398 390788 547634
rect 390440 547366 390788 547398
rect 300952 543454 301300 543486
rect 300952 543218 301008 543454
rect 301244 543218 301300 543454
rect 300952 543134 301300 543218
rect 300952 542898 301008 543134
rect 301244 542898 301300 543134
rect 300952 542866 301300 542898
rect 389760 543454 390108 543486
rect 389760 543218 389816 543454
rect 390052 543218 390108 543454
rect 389760 543134 390108 543218
rect 389760 542898 389816 543134
rect 390052 542898 390108 543134
rect 389760 542866 390108 542898
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 300272 511954 300620 511986
rect 300272 511718 300328 511954
rect 300564 511718 300620 511954
rect 300272 511634 300620 511718
rect 300272 511398 300328 511634
rect 300564 511398 300620 511634
rect 300272 511366 300620 511398
rect 390440 511954 390788 511986
rect 390440 511718 390496 511954
rect 390732 511718 390788 511954
rect 390440 511634 390788 511718
rect 390440 511398 390496 511634
rect 390732 511398 390788 511634
rect 390440 511366 390788 511398
rect 300952 507454 301300 507486
rect 300952 507218 301008 507454
rect 301244 507218 301300 507454
rect 300952 507134 301300 507218
rect 300952 506898 301008 507134
rect 301244 506898 301300 507134
rect 300952 506866 301300 506898
rect 389760 507454 390108 507486
rect 389760 507218 389816 507454
rect 390052 507218 390108 507454
rect 389760 507134 390108 507218
rect 389760 506898 389816 507134
rect 390052 506898 390108 507134
rect 389760 506866 390108 506898
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 312928 489930 312988 490106
rect 312862 489870 312988 489930
rect 314288 489930 314348 490106
rect 315376 489930 315436 490106
rect 317688 489930 317748 490106
rect 314288 489870 314394 489930
rect 315376 489870 315498 489930
rect 312862 487253 312922 489870
rect 314334 488341 314394 489870
rect 314331 488340 314397 488341
rect 314331 488276 314332 488340
rect 314396 488276 314397 488340
rect 314331 488275 314397 488276
rect 315438 488205 315498 489870
rect 317646 489870 317748 489930
rect 318912 489930 318972 490106
rect 320000 489930 320060 490106
rect 321088 489930 321148 490106
rect 322312 489930 322372 490106
rect 323400 489930 323460 490106
rect 318912 489870 318994 489930
rect 320000 489870 320098 489930
rect 321088 489870 321202 489930
rect 315435 488204 315501 488205
rect 315435 488140 315436 488204
rect 315500 488140 315501 488204
rect 315435 488139 315501 488140
rect 317646 487253 317706 489870
rect 318934 487933 318994 489870
rect 318931 487932 318997 487933
rect 318931 487868 318932 487932
rect 318996 487868 318997 487932
rect 318931 487867 318997 487868
rect 320038 487253 320098 489870
rect 321142 487253 321202 489870
rect 322246 489870 322372 489930
rect 323350 489870 323460 489930
rect 324760 489930 324820 490106
rect 325304 489930 325364 490106
rect 325712 489930 325772 490106
rect 330472 489930 330532 490106
rect 335504 489930 335564 490106
rect 324760 489870 324882 489930
rect 325304 489870 325434 489930
rect 325712 489870 325802 489930
rect 330472 489870 330586 489930
rect 322246 487253 322306 489870
rect 323350 487389 323410 489870
rect 323347 487388 323413 487389
rect 323347 487324 323348 487388
rect 323412 487324 323413 487388
rect 323347 487323 323413 487324
rect 324822 487253 324882 489870
rect 325374 489157 325434 489870
rect 325371 489156 325437 489157
rect 325371 489092 325372 489156
rect 325436 489092 325437 489156
rect 325371 489091 325437 489092
rect 325742 487253 325802 489870
rect 330526 488477 330586 489870
rect 335494 489870 335564 489930
rect 340536 489930 340596 490106
rect 345568 489930 345628 490106
rect 350464 489930 350524 490106
rect 340536 489870 340706 489930
rect 345568 489870 345674 489930
rect 335494 488477 335554 489870
rect 340646 488477 340706 489870
rect 345614 488477 345674 489870
rect 350398 489870 350524 489930
rect 355496 489930 355556 490106
rect 360528 489930 360588 490106
rect 355496 489870 355610 489930
rect 350398 488477 350458 489870
rect 355550 488477 355610 489870
rect 360518 489870 360588 489930
rect 360518 488477 360578 489870
rect 330523 488476 330589 488477
rect 330523 488412 330524 488476
rect 330588 488412 330589 488476
rect 330523 488411 330589 488412
rect 335491 488476 335557 488477
rect 335491 488412 335492 488476
rect 335556 488412 335557 488476
rect 335491 488411 335557 488412
rect 340643 488476 340709 488477
rect 340643 488412 340644 488476
rect 340708 488412 340709 488476
rect 340643 488411 340709 488412
rect 345611 488476 345677 488477
rect 345611 488412 345612 488476
rect 345676 488412 345677 488476
rect 345611 488411 345677 488412
rect 350395 488476 350461 488477
rect 350395 488412 350396 488476
rect 350460 488412 350461 488476
rect 350395 488411 350461 488412
rect 355547 488476 355613 488477
rect 355547 488412 355548 488476
rect 355612 488412 355613 488476
rect 355547 488411 355613 488412
rect 360515 488476 360581 488477
rect 360515 488412 360516 488476
rect 360580 488412 360581 488476
rect 360515 488411 360581 488412
rect 312859 487252 312925 487253
rect 312859 487188 312860 487252
rect 312924 487188 312925 487252
rect 312859 487187 312925 487188
rect 317643 487252 317709 487253
rect 317643 487188 317644 487252
rect 317708 487188 317709 487252
rect 317643 487187 317709 487188
rect 320035 487252 320101 487253
rect 320035 487188 320036 487252
rect 320100 487188 320101 487252
rect 320035 487187 320101 487188
rect 321139 487252 321205 487253
rect 321139 487188 321140 487252
rect 321204 487188 321205 487252
rect 321139 487187 321205 487188
rect 322243 487252 322309 487253
rect 322243 487188 322244 487252
rect 322308 487188 322309 487252
rect 322243 487187 322309 487188
rect 324819 487252 324885 487253
rect 324819 487188 324820 487252
rect 324884 487188 324885 487252
rect 324819 487187 324885 487188
rect 325739 487252 325805 487253
rect 325739 487188 325740 487252
rect 325804 487188 325805 487252
rect 325739 487187 325805 487188
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 388794 462454 389414 488000
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 298507 446180 298573 446181
rect 298507 446116 298508 446180
rect 298572 446116 298573 446180
rect 298507 446115 298573 446116
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 298510 19413 298570 446115
rect 319568 439954 319888 439986
rect 319568 439718 319610 439954
rect 319846 439718 319888 439954
rect 319568 439634 319888 439718
rect 319568 439398 319610 439634
rect 319846 439398 319888 439634
rect 319568 439366 319888 439398
rect 350288 439954 350608 439986
rect 350288 439718 350330 439954
rect 350566 439718 350608 439954
rect 350288 439634 350608 439718
rect 350288 439398 350330 439634
rect 350566 439398 350608 439634
rect 350288 439366 350608 439398
rect 381008 439954 381328 439986
rect 381008 439718 381050 439954
rect 381286 439718 381328 439954
rect 381008 439634 381328 439718
rect 381008 439398 381050 439634
rect 381286 439398 381328 439634
rect 381008 439366 381328 439398
rect 304208 435454 304528 435486
rect 304208 435218 304250 435454
rect 304486 435218 304528 435454
rect 304208 435134 304528 435218
rect 304208 434898 304250 435134
rect 304486 434898 304528 435134
rect 304208 434866 304528 434898
rect 334928 435454 335248 435486
rect 334928 435218 334970 435454
rect 335206 435218 335248 435454
rect 334928 435134 335248 435218
rect 334928 434898 334970 435134
rect 335206 434898 335248 435134
rect 334928 434866 335248 434898
rect 365648 435454 365968 435486
rect 365648 435218 365690 435454
rect 365926 435218 365968 435454
rect 365648 435134 365968 435218
rect 365648 434898 365690 435134
rect 365926 434898 365968 435134
rect 365648 434866 365968 434898
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 319568 403954 319888 403986
rect 319568 403718 319610 403954
rect 319846 403718 319888 403954
rect 319568 403634 319888 403718
rect 319568 403398 319610 403634
rect 319846 403398 319888 403634
rect 319568 403366 319888 403398
rect 350288 403954 350608 403986
rect 350288 403718 350330 403954
rect 350566 403718 350608 403954
rect 350288 403634 350608 403718
rect 350288 403398 350330 403634
rect 350566 403398 350608 403634
rect 350288 403366 350608 403398
rect 381008 403954 381328 403986
rect 381008 403718 381050 403954
rect 381286 403718 381328 403954
rect 381008 403634 381328 403718
rect 381008 403398 381050 403634
rect 381286 403398 381328 403634
rect 381008 403366 381328 403398
rect 383331 402932 383397 402933
rect 383331 402868 383332 402932
rect 383396 402868 383397 402932
rect 383331 402867 383397 402868
rect 383334 401573 383394 402867
rect 383331 401572 383397 401573
rect 383331 401508 383332 401572
rect 383396 401508 383397 401572
rect 383331 401507 383397 401508
rect 298794 372454 299414 398000
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298507 19412 298573 19413
rect 298507 19348 298508 19412
rect 298572 19348 298573 19412
rect 298507 19347 298573 19348
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 376954 303914 398000
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 381454 308414 398000
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 385954 312914 398000
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 390454 317414 398000
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 394954 321914 398000
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 367954 330914 398000
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 372454 335414 398000
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 376954 339914 398000
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 385954 348914 398000
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 390454 353414 398000
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 394954 357914 398000
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 363454 362414 398000
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 367954 366914 398000
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 372454 371414 398000
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 376954 375914 398000
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 381454 380414 398000
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 385954 384914 398000
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 691292 411914 700398
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 691292 438914 691398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 691292 443414 695898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 691292 447914 700398
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 691292 474914 691398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 691292 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 691292 483914 700398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 410952 687454 411300 687486
rect 410952 687218 411008 687454
rect 411244 687218 411300 687454
rect 410952 687134 411300 687218
rect 410952 686898 411008 687134
rect 411244 686898 411300 687134
rect 410952 686866 411300 686898
rect 499760 687454 500108 687486
rect 499760 687218 499816 687454
rect 500052 687218 500108 687454
rect 499760 687134 500108 687218
rect 499760 686898 499816 687134
rect 500052 686898 500108 687134
rect 499760 686866 500108 686898
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 410272 655954 410620 655986
rect 410272 655718 410328 655954
rect 410564 655718 410620 655954
rect 410272 655634 410620 655718
rect 410272 655398 410328 655634
rect 410564 655398 410620 655634
rect 410272 655366 410620 655398
rect 500440 655954 500788 655986
rect 500440 655718 500496 655954
rect 500732 655718 500788 655954
rect 500440 655634 500788 655718
rect 500440 655398 500496 655634
rect 500732 655398 500788 655634
rect 500440 655366 500788 655398
rect 410952 651454 411300 651486
rect 410952 651218 411008 651454
rect 411244 651218 411300 651454
rect 410952 651134 411300 651218
rect 410952 650898 411008 651134
rect 411244 650898 411300 651134
rect 410952 650866 411300 650898
rect 499760 651454 500108 651486
rect 499760 651218 499816 651454
rect 500052 651218 500108 651454
rect 499760 651134 500108 651218
rect 499760 650898 499816 651134
rect 500052 650898 500108 651134
rect 499760 650866 500108 650898
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 410272 619954 410620 619986
rect 410272 619718 410328 619954
rect 410564 619718 410620 619954
rect 410272 619634 410620 619718
rect 410272 619398 410328 619634
rect 410564 619398 410620 619634
rect 410272 619366 410620 619398
rect 500440 619954 500788 619986
rect 500440 619718 500496 619954
rect 500732 619718 500788 619954
rect 500440 619634 500788 619718
rect 500440 619398 500496 619634
rect 500732 619398 500788 619634
rect 500440 619366 500788 619398
rect 410952 615454 411300 615486
rect 410952 615218 411008 615454
rect 411244 615218 411300 615454
rect 410952 615134 411300 615218
rect 410952 614898 411008 615134
rect 411244 614898 411300 615134
rect 410952 614866 411300 614898
rect 499760 615454 500108 615486
rect 499760 615218 499816 615454
rect 500052 615218 500108 615454
rect 499760 615134 500108 615218
rect 499760 614898 499816 615134
rect 500052 614898 500108 615134
rect 499760 614866 500108 614898
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 422928 599450 422988 600100
rect 424288 599450 424348 600100
rect 425376 599450 425436 600100
rect 427688 599450 427748 600100
rect 422894 599390 422988 599450
rect 424182 599390 424348 599450
rect 425286 599390 425436 599450
rect 427678 599390 427748 599450
rect 428912 599450 428972 600100
rect 430000 599450 430060 600100
rect 431088 599450 431148 600100
rect 432312 599450 432372 600100
rect 433400 599450 433460 600100
rect 434760 599450 434820 600100
rect 435304 599450 435364 600100
rect 435712 599450 435772 600100
rect 440472 599450 440532 600100
rect 428912 599390 429026 599450
rect 422894 596461 422954 599390
rect 422891 596460 422957 596461
rect 422891 596396 422892 596460
rect 422956 596396 422957 596460
rect 422891 596395 422957 596396
rect 424182 596325 424242 599390
rect 425286 596325 425346 599390
rect 427678 597141 427738 599390
rect 428966 597277 429026 599390
rect 429886 599390 430060 599450
rect 430990 599390 431148 599450
rect 431726 599390 432372 599450
rect 433382 599390 433460 599450
rect 434670 599390 434820 599450
rect 435222 599390 435364 599450
rect 435590 599390 435772 599450
rect 440374 599390 440532 599450
rect 445504 599450 445564 600100
rect 450536 599450 450596 600100
rect 455568 599450 455628 600100
rect 460464 599450 460524 600100
rect 465496 599450 465556 600100
rect 470528 599450 470588 600100
rect 445504 599390 445586 599450
rect 429886 597549 429946 599390
rect 429883 597548 429949 597549
rect 429883 597484 429884 597548
rect 429948 597484 429949 597548
rect 429883 597483 429949 597484
rect 430990 597413 431050 599390
rect 430987 597412 431053 597413
rect 430987 597348 430988 597412
rect 431052 597348 431053 597412
rect 430987 597347 431053 597348
rect 428963 597276 429029 597277
rect 428963 597212 428964 597276
rect 429028 597212 429029 597276
rect 428963 597211 429029 597212
rect 427675 597140 427741 597141
rect 427675 597076 427676 597140
rect 427740 597076 427741 597140
rect 427675 597075 427741 597076
rect 431726 596869 431786 599390
rect 433382 597277 433442 599390
rect 433379 597276 433445 597277
rect 433379 597212 433380 597276
rect 433444 597212 433445 597276
rect 433379 597211 433445 597212
rect 434670 597141 434730 599390
rect 434667 597140 434733 597141
rect 434667 597076 434668 597140
rect 434732 597076 434733 597140
rect 434667 597075 434733 597076
rect 435222 597005 435282 599390
rect 435590 597549 435650 599390
rect 435587 597548 435653 597549
rect 435587 597484 435588 597548
rect 435652 597484 435653 597548
rect 435587 597483 435653 597484
rect 440374 597413 440434 599390
rect 445526 597549 445586 599390
rect 450494 599390 450596 599450
rect 455462 599390 455628 599450
rect 460430 599390 460524 599450
rect 465398 599390 465556 599450
rect 470366 599390 470588 599450
rect 445523 597548 445589 597549
rect 445523 597484 445524 597548
rect 445588 597484 445589 597548
rect 445523 597483 445589 597484
rect 440371 597412 440437 597413
rect 440371 597348 440372 597412
rect 440436 597348 440437 597412
rect 440371 597347 440437 597348
rect 450494 597277 450554 599390
rect 455462 597413 455522 599390
rect 460430 597549 460490 599390
rect 460427 597548 460493 597549
rect 460427 597484 460428 597548
rect 460492 597484 460493 597548
rect 460427 597483 460493 597484
rect 465398 597413 465458 599390
rect 455459 597412 455525 597413
rect 455459 597348 455460 597412
rect 455524 597348 455525 597412
rect 455459 597347 455525 597348
rect 465395 597412 465461 597413
rect 465395 597348 465396 597412
rect 465460 597348 465461 597412
rect 465395 597347 465461 597348
rect 450491 597276 450557 597277
rect 450491 597212 450492 597276
rect 450556 597212 450557 597276
rect 450491 597211 450557 597212
rect 470366 597005 470426 599390
rect 435219 597004 435285 597005
rect 435219 596940 435220 597004
rect 435284 596940 435285 597004
rect 435219 596939 435285 596940
rect 470363 597004 470429 597005
rect 470363 596940 470364 597004
rect 470428 596940 470429 597004
rect 470363 596939 470429 596940
rect 431723 596868 431789 596869
rect 431723 596804 431724 596868
rect 431788 596804 431789 596868
rect 431723 596803 431789 596804
rect 424179 596324 424245 596325
rect 424179 596260 424180 596324
rect 424244 596260 424245 596324
rect 424179 596259 424245 596260
rect 425283 596324 425349 596325
rect 425283 596260 425284 596324
rect 425348 596260 425349 596324
rect 425283 596259 425349 596260
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 410272 547954 410620 547986
rect 410272 547718 410328 547954
rect 410564 547718 410620 547954
rect 410272 547634 410620 547718
rect 410272 547398 410328 547634
rect 410564 547398 410620 547634
rect 410272 547366 410620 547398
rect 500440 547954 500788 547986
rect 500440 547718 500496 547954
rect 500732 547718 500788 547954
rect 500440 547634 500788 547718
rect 500440 547398 500496 547634
rect 500732 547398 500788 547634
rect 500440 547366 500788 547398
rect 410952 543454 411300 543486
rect 410952 543218 411008 543454
rect 411244 543218 411300 543454
rect 410952 543134 411300 543218
rect 410952 542898 411008 543134
rect 411244 542898 411300 543134
rect 410952 542866 411300 542898
rect 499760 543454 500108 543486
rect 499760 543218 499816 543454
rect 500052 543218 500108 543454
rect 499760 543134 500108 543218
rect 499760 542898 499816 543134
rect 500052 542898 500108 543134
rect 499760 542866 500108 542898
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 407803 523700 407869 523701
rect 407803 523636 407804 523700
rect 407868 523636 407869 523700
rect 407803 523635 407869 523636
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 407806 489837 407866 523635
rect 410272 511954 410620 511986
rect 410272 511718 410328 511954
rect 410564 511718 410620 511954
rect 410272 511634 410620 511718
rect 410272 511398 410328 511634
rect 410564 511398 410620 511634
rect 410272 511366 410620 511398
rect 500440 511954 500788 511986
rect 500440 511718 500496 511954
rect 500732 511718 500788 511954
rect 500440 511634 500788 511718
rect 500440 511398 500496 511634
rect 500732 511398 500788 511634
rect 500440 511366 500788 511398
rect 410952 507454 411300 507486
rect 410952 507218 411008 507454
rect 411244 507218 411300 507454
rect 410952 507134 411300 507218
rect 410952 506898 411008 507134
rect 411244 506898 411300 507134
rect 410952 506866 411300 506898
rect 499760 507454 500108 507486
rect 499760 507218 499816 507454
rect 500052 507218 500108 507454
rect 499760 507134 500108 507218
rect 499760 506898 499816 507134
rect 500052 506898 500108 507134
rect 499760 506866 500108 506898
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 422928 489930 422988 490106
rect 424288 489930 424348 490106
rect 425376 489930 425436 490106
rect 427688 489930 427748 490106
rect 422894 489870 422988 489930
rect 424182 489870 424348 489930
rect 425286 489870 425436 489930
rect 427678 489870 427748 489930
rect 428912 489930 428972 490106
rect 430000 489930 430060 490106
rect 431088 489930 431148 490106
rect 432312 489930 432372 490106
rect 433400 489930 433460 490106
rect 428912 489870 429026 489930
rect 407803 489836 407869 489837
rect 407803 489772 407804 489836
rect 407868 489772 407869 489836
rect 407803 489771 407869 489772
rect 422894 488477 422954 489870
rect 424182 488477 424242 489870
rect 422891 488476 422957 488477
rect 422891 488412 422892 488476
rect 422956 488412 422957 488476
rect 422891 488411 422957 488412
rect 424179 488476 424245 488477
rect 424179 488412 424180 488476
rect 424244 488412 424245 488476
rect 424179 488411 424245 488412
rect 425286 488341 425346 489870
rect 425283 488340 425349 488341
rect 425283 488276 425284 488340
rect 425348 488276 425349 488340
rect 425283 488275 425349 488276
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 484954 411914 488000
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 453454 416414 488000
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 457954 420914 488000
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 462454 425414 488000
rect 427678 487797 427738 489870
rect 428966 488205 429026 489870
rect 429886 489870 430060 489930
rect 430990 489870 431148 489930
rect 432278 489870 432372 489930
rect 433382 489870 433460 489930
rect 434760 489930 434820 490106
rect 435304 489930 435364 490106
rect 435712 489930 435772 490106
rect 440472 489930 440532 490106
rect 434760 489870 434914 489930
rect 429886 488205 429946 489870
rect 430990 488341 431050 489870
rect 430987 488340 431053 488341
rect 430987 488276 430988 488340
rect 431052 488276 431053 488340
rect 430987 488275 431053 488276
rect 428963 488204 429029 488205
rect 428963 488140 428964 488204
rect 429028 488140 429029 488204
rect 428963 488139 429029 488140
rect 429883 488204 429949 488205
rect 429883 488140 429884 488204
rect 429948 488140 429949 488204
rect 429883 488139 429949 488140
rect 427675 487796 427741 487797
rect 427675 487732 427676 487796
rect 427740 487732 427741 487796
rect 427675 487731 427741 487732
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 466954 429914 488000
rect 432278 487661 432338 489870
rect 432275 487660 432341 487661
rect 432275 487596 432276 487660
rect 432340 487596 432341 487660
rect 432275 487595 432341 487596
rect 433382 487389 433442 489870
rect 433379 487388 433445 487389
rect 433379 487324 433380 487388
rect 433444 487324 433445 487388
rect 433379 487323 433445 487324
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 471454 434414 488000
rect 434854 487253 434914 489870
rect 435222 489870 435364 489930
rect 435590 489870 435772 489930
rect 440374 489870 440532 489930
rect 445504 489930 445564 490106
rect 450536 489930 450596 490106
rect 455568 489930 455628 490106
rect 460464 489930 460524 490106
rect 465496 489930 465556 490106
rect 445504 489870 445586 489930
rect 435222 488477 435282 489870
rect 435219 488476 435285 488477
rect 435219 488412 435220 488476
rect 435284 488412 435285 488476
rect 435219 488411 435285 488412
rect 435590 488205 435650 489870
rect 440374 488477 440434 489870
rect 445526 488477 445586 489870
rect 450494 489870 450596 489930
rect 455462 489870 455628 489930
rect 460430 489870 460524 489930
rect 465398 489870 465556 489930
rect 470528 489930 470588 490106
rect 470528 489870 470794 489930
rect 450494 488477 450554 489870
rect 440371 488476 440437 488477
rect 440371 488412 440372 488476
rect 440436 488412 440437 488476
rect 440371 488411 440437 488412
rect 445523 488476 445589 488477
rect 445523 488412 445524 488476
rect 445588 488412 445589 488476
rect 445523 488411 445589 488412
rect 450491 488476 450557 488477
rect 450491 488412 450492 488476
rect 450556 488412 450557 488476
rect 450491 488411 450557 488412
rect 435587 488204 435653 488205
rect 435587 488140 435588 488204
rect 435652 488140 435653 488204
rect 435587 488139 435653 488140
rect 455462 488069 455522 489870
rect 455459 488068 455525 488069
rect 455459 488004 455460 488068
rect 455524 488004 455525 488068
rect 455459 488003 455525 488004
rect 434851 487252 434917 487253
rect 434851 487188 434852 487252
rect 434916 487188 434917 487252
rect 434851 487187 434917 487188
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 475954 438914 488000
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 480454 443414 488000
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 484954 447914 488000
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 453454 452414 488000
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 457954 456914 488000
rect 460430 487933 460490 489870
rect 465398 488341 465458 489870
rect 465395 488340 465461 488341
rect 465395 488276 465396 488340
rect 465460 488276 465461 488340
rect 465395 488275 465461 488276
rect 470734 488069 470794 489870
rect 470731 488068 470797 488069
rect 470731 488004 470732 488068
rect 470796 488004 470797 488068
rect 470731 488003 470797 488004
rect 460427 487932 460493 487933
rect 460427 487868 460428 487932
rect 460492 487868 460493 487932
rect 460427 487867 460493 487868
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 462454 461414 488000
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 466954 465914 488000
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 471454 470414 488000
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 475954 474914 488000
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 480454 479414 488000
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 484954 483914 488000
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 453454 488414 488000
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 457954 492914 488000
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 462454 497414 488000
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 466954 501914 488000
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 81008 687218 81244 687454
rect 81008 686898 81244 687134
rect 169816 687218 170052 687454
rect 169816 686898 170052 687134
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 80328 655718 80564 655954
rect 80328 655398 80564 655634
rect 170496 655718 170732 655954
rect 170496 655398 170732 655634
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 81008 651218 81244 651454
rect 81008 650898 81244 651134
rect 169816 651218 170052 651454
rect 169816 650898 170052 651134
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 80328 619718 80564 619954
rect 80328 619398 80564 619634
rect 170496 619718 170732 619954
rect 170496 619398 170732 619634
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 81008 615218 81244 615454
rect 81008 614898 81244 615134
rect 169816 615218 170052 615454
rect 169816 614898 170052 615134
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 80328 547718 80564 547954
rect 80328 547398 80564 547634
rect 170496 547718 170732 547954
rect 170496 547398 170732 547634
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 81008 543218 81244 543454
rect 81008 542898 81244 543134
rect 169816 543218 170052 543454
rect 169816 542898 170052 543134
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 80328 511718 80564 511954
rect 80328 511398 80564 511634
rect 170496 511718 170732 511954
rect 170496 511398 170732 511634
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 81008 507218 81244 507454
rect 81008 506898 81244 507134
rect 169816 507218 170052 507454
rect 169816 506898 170052 507134
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 191008 687218 191244 687454
rect 191008 686898 191244 687134
rect 279816 687218 280052 687454
rect 279816 686898 280052 687134
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 190328 655718 190564 655954
rect 190328 655398 190564 655634
rect 280496 655718 280732 655954
rect 280496 655398 280732 655634
rect 191008 651218 191244 651454
rect 191008 650898 191244 651134
rect 279816 651218 280052 651454
rect 279816 650898 280052 651134
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190328 619718 190564 619954
rect 190328 619398 190564 619634
rect 280496 619718 280732 619954
rect 280496 619398 280732 619634
rect 191008 615218 191244 615454
rect 191008 614898 191244 615134
rect 279816 615218 280052 615454
rect 279816 614898 280052 615134
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 190328 547718 190564 547954
rect 190328 547398 190564 547634
rect 280496 547718 280732 547954
rect 280496 547398 280732 547634
rect 191008 543218 191244 543454
rect 191008 542898 191244 543134
rect 279816 543218 280052 543454
rect 279816 542898 280052 543134
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 190328 511718 190564 511954
rect 190328 511398 190564 511634
rect 280496 511718 280732 511954
rect 280496 511398 280732 511634
rect 191008 507218 191244 507454
rect 191008 506898 191244 507134
rect 279816 507218 280052 507454
rect 279816 506898 280052 507134
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 219610 439718 219846 439954
rect 219610 439398 219846 439634
rect 250330 439718 250566 439954
rect 250330 439398 250566 439634
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 219610 403718 219846 403954
rect 219610 403398 219846 403634
rect 250330 403718 250566 403954
rect 250330 403398 250566 403634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 301008 687218 301244 687454
rect 301008 686898 301244 687134
rect 389816 687218 390052 687454
rect 389816 686898 390052 687134
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 300328 655718 300564 655954
rect 300328 655398 300564 655634
rect 390496 655718 390732 655954
rect 390496 655398 390732 655634
rect 301008 651218 301244 651454
rect 301008 650898 301244 651134
rect 389816 651218 390052 651454
rect 389816 650898 390052 651134
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 300328 619718 300564 619954
rect 300328 619398 300564 619634
rect 390496 619718 390732 619954
rect 390496 619398 390732 619634
rect 301008 615218 301244 615454
rect 301008 614898 301244 615134
rect 389816 615218 390052 615454
rect 389816 614898 390052 615134
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 300328 547718 300564 547954
rect 300328 547398 300564 547634
rect 390496 547718 390732 547954
rect 390496 547398 390732 547634
rect 301008 543218 301244 543454
rect 301008 542898 301244 543134
rect 389816 543218 390052 543454
rect 389816 542898 390052 543134
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 300328 511718 300564 511954
rect 300328 511398 300564 511634
rect 390496 511718 390732 511954
rect 390496 511398 390732 511634
rect 301008 507218 301244 507454
rect 301008 506898 301244 507134
rect 389816 507218 390052 507454
rect 389816 506898 390052 507134
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 319610 439718 319846 439954
rect 319610 439398 319846 439634
rect 350330 439718 350566 439954
rect 350330 439398 350566 439634
rect 381050 439718 381286 439954
rect 381050 439398 381286 439634
rect 304250 435218 304486 435454
rect 304250 434898 304486 435134
rect 334970 435218 335206 435454
rect 334970 434898 335206 435134
rect 365690 435218 365926 435454
rect 365690 434898 365926 435134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 319610 403718 319846 403954
rect 319610 403398 319846 403634
rect 350330 403718 350566 403954
rect 350330 403398 350566 403634
rect 381050 403718 381286 403954
rect 381050 403398 381286 403634
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 411008 687218 411244 687454
rect 411008 686898 411244 687134
rect 499816 687218 500052 687454
rect 499816 686898 500052 687134
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 410328 655718 410564 655954
rect 410328 655398 410564 655634
rect 500496 655718 500732 655954
rect 500496 655398 500732 655634
rect 411008 651218 411244 651454
rect 411008 650898 411244 651134
rect 499816 651218 500052 651454
rect 499816 650898 500052 651134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 410328 619718 410564 619954
rect 410328 619398 410564 619634
rect 500496 619718 500732 619954
rect 500496 619398 500732 619634
rect 411008 615218 411244 615454
rect 411008 614898 411244 615134
rect 499816 615218 500052 615454
rect 499816 614898 500052 615134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 410328 547718 410564 547954
rect 410328 547398 410564 547634
rect 500496 547718 500732 547954
rect 500496 547398 500732 547634
rect 411008 543218 411244 543454
rect 411008 542898 411244 543134
rect 499816 543218 500052 543454
rect 499816 542898 500052 543134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 410328 511718 410564 511954
rect 410328 511398 410564 511634
rect 500496 511718 500732 511954
rect 500496 511398 500732 511634
rect 411008 507218 411244 507454
rect 411008 506898 411244 507134
rect 499816 507218 500052 507454
rect 499816 506898 500052 507134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 81008 687454
rect 81244 687218 169816 687454
rect 170052 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 191008 687454
rect 191244 687218 279816 687454
rect 280052 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 301008 687454
rect 301244 687218 389816 687454
rect 390052 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 411008 687454
rect 411244 687218 499816 687454
rect 500052 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 81008 687134
rect 81244 686898 169816 687134
rect 170052 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 191008 687134
rect 191244 686898 279816 687134
rect 280052 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 301008 687134
rect 301244 686898 389816 687134
rect 390052 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 411008 687134
rect 411244 686898 499816 687134
rect 500052 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 80328 655954
rect 80564 655718 170496 655954
rect 170732 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 190328 655954
rect 190564 655718 280496 655954
rect 280732 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 300328 655954
rect 300564 655718 390496 655954
rect 390732 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 410328 655954
rect 410564 655718 500496 655954
rect 500732 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 80328 655634
rect 80564 655398 170496 655634
rect 170732 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 190328 655634
rect 190564 655398 280496 655634
rect 280732 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 300328 655634
rect 300564 655398 390496 655634
rect 390732 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 410328 655634
rect 410564 655398 500496 655634
rect 500732 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 81008 651454
rect 81244 651218 169816 651454
rect 170052 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 191008 651454
rect 191244 651218 279816 651454
rect 280052 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 301008 651454
rect 301244 651218 389816 651454
rect 390052 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 411008 651454
rect 411244 651218 499816 651454
rect 500052 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 81008 651134
rect 81244 650898 169816 651134
rect 170052 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 191008 651134
rect 191244 650898 279816 651134
rect 280052 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 301008 651134
rect 301244 650898 389816 651134
rect 390052 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 411008 651134
rect 411244 650898 499816 651134
rect 500052 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 80328 619954
rect 80564 619718 170496 619954
rect 170732 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 190328 619954
rect 190564 619718 280496 619954
rect 280732 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 300328 619954
rect 300564 619718 390496 619954
rect 390732 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 410328 619954
rect 410564 619718 500496 619954
rect 500732 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 80328 619634
rect 80564 619398 170496 619634
rect 170732 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 190328 619634
rect 190564 619398 280496 619634
rect 280732 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 300328 619634
rect 300564 619398 390496 619634
rect 390732 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 410328 619634
rect 410564 619398 500496 619634
rect 500732 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 81008 615454
rect 81244 615218 169816 615454
rect 170052 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 191008 615454
rect 191244 615218 279816 615454
rect 280052 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 301008 615454
rect 301244 615218 389816 615454
rect 390052 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 411008 615454
rect 411244 615218 499816 615454
rect 500052 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 81008 615134
rect 81244 614898 169816 615134
rect 170052 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 191008 615134
rect 191244 614898 279816 615134
rect 280052 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 301008 615134
rect 301244 614898 389816 615134
rect 390052 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 411008 615134
rect 411244 614898 499816 615134
rect 500052 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 80328 547954
rect 80564 547718 170496 547954
rect 170732 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 190328 547954
rect 190564 547718 280496 547954
rect 280732 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 300328 547954
rect 300564 547718 390496 547954
rect 390732 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 410328 547954
rect 410564 547718 500496 547954
rect 500732 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 80328 547634
rect 80564 547398 170496 547634
rect 170732 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 190328 547634
rect 190564 547398 280496 547634
rect 280732 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 300328 547634
rect 300564 547398 390496 547634
rect 390732 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 410328 547634
rect 410564 547398 500496 547634
rect 500732 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 81008 543454
rect 81244 543218 169816 543454
rect 170052 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 191008 543454
rect 191244 543218 279816 543454
rect 280052 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 301008 543454
rect 301244 543218 389816 543454
rect 390052 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 411008 543454
rect 411244 543218 499816 543454
rect 500052 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 81008 543134
rect 81244 542898 169816 543134
rect 170052 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 191008 543134
rect 191244 542898 279816 543134
rect 280052 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 301008 543134
rect 301244 542898 389816 543134
rect 390052 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 411008 543134
rect 411244 542898 499816 543134
rect 500052 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 80328 511954
rect 80564 511718 170496 511954
rect 170732 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 190328 511954
rect 190564 511718 280496 511954
rect 280732 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 300328 511954
rect 300564 511718 390496 511954
rect 390732 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 410328 511954
rect 410564 511718 500496 511954
rect 500732 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 80328 511634
rect 80564 511398 170496 511634
rect 170732 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 190328 511634
rect 190564 511398 280496 511634
rect 280732 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 300328 511634
rect 300564 511398 390496 511634
rect 390732 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 410328 511634
rect 410564 511398 500496 511634
rect 500732 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 81008 507454
rect 81244 507218 169816 507454
rect 170052 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 191008 507454
rect 191244 507218 279816 507454
rect 280052 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 301008 507454
rect 301244 507218 389816 507454
rect 390052 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 411008 507454
rect 411244 507218 499816 507454
rect 500052 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 81008 507134
rect 81244 506898 169816 507134
rect 170052 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 191008 507134
rect 191244 506898 279816 507134
rect 280052 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 301008 507134
rect 301244 506898 389816 507134
rect 390052 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 411008 507134
rect 411244 506898 499816 507134
rect 500052 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 219610 439954
rect 219846 439718 250330 439954
rect 250566 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 319610 439954
rect 319846 439718 350330 439954
rect 350566 439718 381050 439954
rect 381286 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 219610 439634
rect 219846 439398 250330 439634
rect 250566 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 319610 439634
rect 319846 439398 350330 439634
rect 350566 439398 381050 439634
rect 381286 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 304250 435454
rect 304486 435218 334970 435454
rect 335206 435218 365690 435454
rect 365926 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 304250 435134
rect 304486 434898 334970 435134
rect 335206 434898 365690 435134
rect 365926 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 219610 403954
rect 219846 403718 250330 403954
rect 250566 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 319610 403954
rect 319846 403718 350330 403954
rect 350566 403718 381050 403954
rect 381286 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 219610 403634
rect 219846 403398 250330 403634
rect 250566 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 319610 403634
rect 319846 403398 350330 403634
rect 350566 403398 381050 403634
rect 381286 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use cpu  cpu0
timestamp 0
transform 1 0 300000 0 1 400000
box 0 0 84000 56000
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword0
timestamp 0
transform 1 0 80000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword1
timestamp 0
transform 1 0 190000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword2
timestamp 0
transform 1 0 300000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword3
timestamp 0
transform 1 0 410000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword0
timestamp 0
transform 1 0 80000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword1
timestamp 0
transform 1 0 190000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword2
timestamp 0
transform 1 0 300000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword3
timestamp 0
transform 1 0 410000 0 1 490000
box 0 0 91060 89292
use soc_config  mprj
timestamp 0
transform 1 0 200000 0 1 400000
box 1066 0 64898 44000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 691292 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 691292 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 691292 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 691292 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 691292 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 691292 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 691292 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 691292 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 691292 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 691292 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 691292 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 691292 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 691292 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 691292 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 691292 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 691292 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 691292 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 691292 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 691292 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 691292 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 691292 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 691292 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 691292 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 691292 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 446000 231914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 691292 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 446000 267914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 691292 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 691292 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 691292 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 691292 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 691292 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 691292 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 691292 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
