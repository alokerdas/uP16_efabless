magic
tech sky130B
magscale 1 2
timestamp 1669281156
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 404998 700544 405004 700596
rect 405056 700584 405062 700596
rect 413646 700584 413652 700596
rect 405056 700556 413652 700584
rect 405056 700544 405062 700556
rect 413646 700544 413652 700556
rect 413704 700544 413710 700596
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 182818 700516 182824 700528
rect 154172 700488 182824 700516
rect 154172 700476 154178 700488
rect 182818 700476 182824 700488
rect 182876 700476 182882 700528
rect 296070 700476 296076 700528
rect 296128 700516 296134 700528
rect 300118 700516 300124 700528
rect 296128 700488 300124 700516
rect 296128 700476 296134 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 409138 700476 409144 700528
rect 409196 700516 409202 700528
rect 429838 700516 429844 700528
rect 409196 700488 429844 700516
rect 409196 700476 409202 700488
rect 429838 700476 429844 700488
rect 429896 700476 429902 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 178678 700448 178684 700460
rect 137888 700420 178684 700448
rect 137888 700408 137894 700420
rect 178678 700408 178684 700420
rect 178736 700408 178742 700460
rect 188890 700408 188896 700460
rect 188948 700448 188954 700460
rect 202782 700448 202788 700460
rect 188948 700420 202788 700448
rect 188948 700408 188954 700420
rect 202782 700408 202788 700420
rect 202840 700408 202846 700460
rect 293218 700408 293224 700460
rect 293276 700448 293282 700460
rect 332502 700448 332508 700460
rect 293276 700420 332508 700448
rect 293276 700408 293282 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 403618 700408 403624 700460
rect 403676 700448 403682 700460
rect 462314 700448 462320 700460
rect 403676 700420 462320 700448
rect 403676 700408 403682 700420
rect 462314 700408 462320 700420
rect 462372 700408 462378 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 174538 700380 174544 700392
rect 105504 700352 174544 700380
rect 105504 700340 105510 700352
rect 174538 700340 174544 700352
rect 174596 700340 174602 700392
rect 188982 700340 188988 700392
rect 189040 700380 189046 700392
rect 218974 700380 218980 700392
rect 189040 700352 218980 700380
rect 189040 700340 189046 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 291838 700340 291844 700392
rect 291896 700380 291902 700392
rect 348786 700380 348792 700392
rect 291896 700352 348792 700380
rect 291896 700340 291902 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 399478 700340 399484 700392
rect 399536 700380 399542 700392
rect 478506 700380 478512 700392
rect 399536 700352 478512 700380
rect 399536 700340 399542 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 184198 700312 184204 700324
rect 89220 700284 184204 700312
rect 89220 700272 89226 700284
rect 184198 700272 184204 700284
rect 184256 700272 184262 700324
rect 188798 700272 188804 700324
rect 188856 700312 188862 700324
rect 235166 700312 235172 700324
rect 188856 700284 235172 700312
rect 188856 700272 188862 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 281534 700312 281540 700324
rect 267700 700284 281540 700312
rect 267700 700272 267706 700284
rect 281534 700272 281540 700284
rect 281592 700272 281598 700324
rect 295978 700272 295984 700324
rect 296036 700312 296042 700324
rect 364978 700312 364984 700324
rect 296036 700284 364984 700312
rect 296036 700272 296042 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 406378 700272 406384 700324
rect 406436 700312 406442 700324
rect 494790 700312 494796 700324
rect 406436 700284 494796 700312
rect 406436 700272 406442 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 509878 700272 509884 700324
rect 509936 700312 509942 700324
rect 559650 700312 559656 700324
rect 509936 700284 559656 700312
rect 509936 700272 509942 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171778 699700 171784 699712
rect 170364 699672 171784 699700
rect 170364 699660 170370 699672
rect 171778 699660 171784 699672
rect 171836 699660 171842 699712
rect 395338 699660 395344 699712
rect 395396 699700 395402 699712
rect 397454 699700 397460 699712
rect 395396 699672 397460 699700
rect 395396 699660 395402 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 286318 696940 286324 696992
rect 286376 696980 286382 696992
rect 580166 696980 580172 696992
rect 286376 696952 580172 696980
rect 286376 696940 286382 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 508498 670692 508504 670744
rect 508556 670732 508562 670744
rect 580166 670732 580172 670744
rect 508556 670704 580172 670732
rect 508556 670692 508562 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 512638 643084 512644 643136
rect 512696 643124 512702 643136
rect 580166 643124 580172 643136
rect 512696 643096 580172 643124
rect 512696 643084 512702 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 501598 630640 501604 630692
rect 501656 630680 501662 630692
rect 579982 630680 579988 630692
rect 501656 630652 579988 630680
rect 501656 630640 501662 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 504358 616836 504364 616888
rect 504416 616876 504422 616888
rect 580166 616876 580172 616888
rect 504416 616848 580172 616876
rect 504416 616836 504422 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 297358 600244 297364 600296
rect 297416 600284 297422 600296
rect 297818 600284 297824 600296
rect 297416 600256 297824 600284
rect 297416 600244 297422 600256
rect 297818 600244 297824 600256
rect 297876 600244 297882 600296
rect 78122 599972 78128 600024
rect 78180 600012 78186 600024
rect 187234 600012 187240 600024
rect 78180 599984 187240 600012
rect 78180 599972 78186 599984
rect 187234 599972 187240 599984
rect 187292 599972 187298 600024
rect 297818 599972 297824 600024
rect 297876 600012 297882 600024
rect 408034 600012 408040 600024
rect 297876 599984 408040 600012
rect 297876 599972 297882 599984
rect 408034 599972 408040 599984
rect 408092 599972 408098 600024
rect 78030 599904 78036 599956
rect 78088 599944 78094 599956
rect 187142 599944 187148 599956
rect 78088 599916 187148 599944
rect 78088 599904 78094 599916
rect 187142 599904 187148 599916
rect 187200 599904 187206 599956
rect 78582 599836 78588 599888
rect 78640 599876 78646 599888
rect 187326 599876 187332 599888
rect 78640 599848 187332 599876
rect 78640 599836 78646 599848
rect 187326 599836 187332 599848
rect 187384 599836 187390 599888
rect 78214 599768 78220 599820
rect 78272 599808 78278 599820
rect 186866 599808 186872 599820
rect 78272 599780 186872 599808
rect 78272 599768 78278 599780
rect 186866 599768 186872 599780
rect 186924 599768 186930 599820
rect 78398 599700 78404 599752
rect 78456 599740 78462 599752
rect 187050 599740 187056 599752
rect 78456 599712 187056 599740
rect 78456 599700 78462 599712
rect 187050 599700 187056 599712
rect 187108 599700 187114 599752
rect 78490 599632 78496 599684
rect 78548 599672 78554 599684
rect 186958 599672 186964 599684
rect 78548 599644 186964 599672
rect 78548 599632 78554 599644
rect 186958 599632 186964 599644
rect 187016 599632 187022 599684
rect 297910 598884 297916 598936
rect 297968 598924 297974 598936
rect 407942 598924 407948 598936
rect 297968 598896 407948 598924
rect 297968 598884 297974 598896
rect 407942 598884 407948 598896
rect 408000 598884 408006 598936
rect 297450 598816 297456 598868
rect 297508 598856 297514 598868
rect 408126 598856 408132 598868
rect 297508 598828 408132 598856
rect 297508 598816 297514 598828
rect 408126 598816 408132 598828
rect 408184 598816 408190 598868
rect 297542 598748 297548 598800
rect 297600 598788 297606 598800
rect 407574 598788 407580 598800
rect 297600 598760 407580 598788
rect 297600 598748 297606 598760
rect 407574 598748 407580 598760
rect 407632 598748 407638 598800
rect 297266 598000 297272 598052
rect 297324 598040 297330 598052
rect 297910 598040 297916 598052
rect 297324 598012 297916 598040
rect 297324 598000 297330 598012
rect 297910 598000 297916 598012
rect 297968 598000 297974 598052
rect 102870 597252 102876 597304
rect 102928 597292 102934 597304
rect 212442 597292 212448 597304
rect 102928 597264 212448 597292
rect 102928 597252 102934 597264
rect 212442 597252 212448 597264
rect 212500 597252 212506 597304
rect 284294 597252 284300 597304
rect 284352 597292 284358 597304
rect 325786 597292 325792 597304
rect 284352 597264 325792 597292
rect 284352 597252 284358 597264
rect 325786 597252 325792 597264
rect 325844 597292 325850 597304
rect 434714 597292 434720 597304
rect 325844 597264 434720 597292
rect 325844 597252 325850 597264
rect 434714 597252 434720 597264
rect 434772 597252 434778 597304
rect 106090 597184 106096 597236
rect 106148 597224 106154 597236
rect 215938 597224 215944 597236
rect 106148 597196 215944 597224
rect 106148 597184 106154 597196
rect 215938 597184 215944 597196
rect 215996 597184 216002 597236
rect 319438 597184 319444 597236
rect 319496 597224 319502 597236
rect 427814 597224 427820 597236
rect 319496 597196 427820 597224
rect 319496 597184 319502 597196
rect 427814 597184 427820 597196
rect 427872 597184 427878 597236
rect 103422 597116 103428 597168
rect 103480 597156 103486 597168
rect 213822 597156 213828 597168
rect 103480 597128 213828 597156
rect 103480 597116 103486 597128
rect 213822 597116 213828 597128
rect 213880 597116 213886 597168
rect 318334 597116 318340 597168
rect 318392 597156 318398 597168
rect 426434 597156 426440 597168
rect 318392 597128 426440 597156
rect 318392 597116 318398 597128
rect 426434 597116 426440 597128
rect 426492 597116 426498 597168
rect 104802 597048 104808 597100
rect 104860 597088 104866 597100
rect 214834 597088 214840 597100
rect 104860 597060 214840 597088
rect 104860 597048 104866 597060
rect 214834 597048 214840 597060
rect 214892 597048 214898 597100
rect 319254 597048 319260 597100
rect 319312 597088 319318 597100
rect 320082 597088 320088 597100
rect 319312 597060 320088 597088
rect 319312 597048 319318 597060
rect 320082 597048 320088 597060
rect 320140 597088 320146 597100
rect 429194 597088 429200 597100
rect 320140 597060 429200 597088
rect 320140 597048 320146 597060
rect 429194 597048 429200 597060
rect 429252 597048 429258 597100
rect 100662 596980 100668 597032
rect 100720 597020 100726 597032
rect 210050 597020 210056 597032
rect 100720 596992 210056 597020
rect 100720 596980 100726 596992
rect 210050 596980 210056 596992
rect 210108 597020 210114 597032
rect 211062 597020 211068 597032
rect 210108 596992 211068 597020
rect 210108 596980 210114 596992
rect 211062 596980 211068 596992
rect 211120 596980 211126 597032
rect 320910 596980 320916 597032
rect 320968 597020 320974 597032
rect 430574 597020 430580 597032
rect 320968 596992 430580 597020
rect 320968 596980 320974 596992
rect 430574 596980 430580 596992
rect 430632 596980 430638 597032
rect 97902 596912 97908 596964
rect 97960 596952 97966 596964
rect 207106 596952 207112 596964
rect 97960 596924 207112 596952
rect 97960 596912 97966 596924
rect 207106 596912 207112 596924
rect 207164 596912 207170 596964
rect 324406 596912 324412 596964
rect 324464 596952 324470 596964
rect 434714 596952 434720 596964
rect 324464 596924 434720 596952
rect 324464 596912 324470 596924
rect 434714 596912 434720 596924
rect 434772 596912 434778 596964
rect 99282 596844 99288 596896
rect 99340 596884 99346 596896
rect 208394 596884 208400 596896
rect 99340 596856 208400 596884
rect 99340 596844 99346 596856
rect 208394 596844 208400 596856
rect 208452 596844 208458 596896
rect 212442 596844 212448 596896
rect 212500 596884 212506 596896
rect 284570 596884 284576 596896
rect 212500 596856 284576 596884
rect 212500 596844 212506 596856
rect 284570 596844 284576 596856
rect 284628 596844 284634 596896
rect 321554 596844 321560 596896
rect 321612 596884 321618 596896
rect 322290 596884 322296 596896
rect 321612 596856 322296 596884
rect 321612 596844 321618 596856
rect 322290 596844 322296 596856
rect 322348 596884 322354 596896
rect 431954 596884 431960 596896
rect 322348 596856 431960 596884
rect 322348 596844 322354 596856
rect 431954 596844 431960 596856
rect 432012 596844 432018 596896
rect 102042 596776 102048 596828
rect 102100 596816 102106 596828
rect 102100 596788 200114 596816
rect 102100 596776 102106 596788
rect 140682 596504 140688 596556
rect 140740 596544 140746 596556
rect 172238 596544 172244 596556
rect 140740 596516 172244 596544
rect 140740 596504 140746 596516
rect 172238 596504 172244 596516
rect 172296 596504 172302 596556
rect 200086 596544 200114 596788
rect 214834 596776 214840 596828
rect 214892 596816 214898 596828
rect 284386 596816 284392 596828
rect 214892 596788 284392 596816
rect 214892 596776 214898 596788
rect 284386 596776 284392 596788
rect 284444 596776 284450 596828
rect 299198 596776 299204 596828
rect 299256 596816 299262 596828
rect 313274 596816 313280 596828
rect 299256 596788 313280 596816
rect 299256 596776 299262 596788
rect 313274 596776 313280 596788
rect 313332 596776 313338 596828
rect 322934 596776 322940 596828
rect 322992 596816 322998 596828
rect 433334 596816 433340 596828
rect 322992 596788 433340 596816
rect 322992 596776 322998 596788
rect 433334 596776 433340 596788
rect 433392 596776 433398 596828
rect 280982 596708 280988 596760
rect 281040 596748 281046 596760
rect 318334 596748 318340 596760
rect 281040 596720 318340 596748
rect 281040 596708 281046 596720
rect 318334 596708 318340 596720
rect 318392 596708 318398 596760
rect 215938 596640 215944 596692
rect 215996 596680 216002 596692
rect 284294 596680 284300 596692
rect 215996 596652 284300 596680
rect 215996 596640 216002 596652
rect 284294 596640 284300 596652
rect 284352 596640 284358 596692
rect 299290 596640 299296 596692
rect 299348 596680 299354 596692
rect 314654 596680 314660 596692
rect 299348 596652 314660 596680
rect 299348 596640 299354 596652
rect 314654 596640 314660 596652
rect 314712 596640 314718 596692
rect 283098 596572 283104 596624
rect 283156 596612 283162 596624
rect 319254 596612 319260 596624
rect 283156 596584 319260 596612
rect 283156 596572 283162 596584
rect 319254 596572 319260 596584
rect 319312 596572 319318 596624
rect 211154 596544 211160 596556
rect 200086 596516 211160 596544
rect 211154 596504 211160 596516
rect 211212 596544 211218 596556
rect 283006 596544 283012 596556
rect 211212 596516 283012 596544
rect 211212 596504 211218 596516
rect 283006 596504 283012 596516
rect 283064 596544 283070 596556
rect 320910 596544 320916 596556
rect 283064 596516 320916 596544
rect 283064 596504 283070 596516
rect 320910 596504 320916 596516
rect 320968 596504 320974 596556
rect 408126 596504 408132 596556
rect 408184 596544 408190 596556
rect 422570 596544 422576 596556
rect 408184 596516 422576 596544
rect 408184 596504 408190 596516
rect 422570 596504 422576 596516
rect 422628 596504 422634 596556
rect 136542 596436 136548 596488
rect 136600 596476 136606 596488
rect 173342 596476 173348 596488
rect 136600 596448 173348 596476
rect 136600 596436 136606 596448
rect 173342 596436 173348 596448
rect 173400 596436 173406 596488
rect 213822 596436 213828 596488
rect 213880 596476 213886 596488
rect 284478 596476 284484 596488
rect 213880 596448 284484 596476
rect 213880 596436 213886 596448
rect 284478 596436 284484 596448
rect 284536 596436 284542 596488
rect 284570 596436 284576 596488
rect 284628 596476 284634 596488
rect 321554 596476 321560 596488
rect 284628 596448 321560 596476
rect 284628 596436 284634 596448
rect 321554 596436 321560 596448
rect 321612 596436 321618 596488
rect 408034 596436 408040 596488
rect 408092 596476 408098 596488
rect 423674 596476 423680 596488
rect 408092 596448 423680 596476
rect 408092 596436 408098 596448
rect 423674 596436 423680 596448
rect 423732 596436 423738 596488
rect 131022 596368 131028 596420
rect 131080 596408 131086 596420
rect 171870 596408 171876 596420
rect 131080 596380 171876 596408
rect 131080 596368 131086 596380
rect 171870 596368 171876 596380
rect 171928 596368 171934 596420
rect 208394 596368 208400 596420
rect 208452 596408 208458 596420
rect 281626 596408 281632 596420
rect 208452 596380 281632 596408
rect 208452 596368 208458 596380
rect 281626 596368 281632 596380
rect 281684 596408 281690 596420
rect 319438 596408 319444 596420
rect 281684 596380 319444 596408
rect 281684 596368 281690 596380
rect 319438 596368 319444 596380
rect 319496 596368 319502 596420
rect 407942 596368 407948 596420
rect 408000 596408 408006 596420
rect 425054 596408 425060 596420
rect 408000 596380 425060 596408
rect 408000 596368 408006 596380
rect 425054 596368 425060 596380
rect 425112 596368 425118 596420
rect 79870 596300 79876 596352
rect 79928 596340 79934 596352
rect 92474 596340 92480 596352
rect 79928 596312 92480 596340
rect 79928 596300 79934 596312
rect 92474 596300 92480 596312
rect 92532 596300 92538 596352
rect 126882 596300 126888 596352
rect 126940 596340 126946 596352
rect 173158 596340 173164 596352
rect 126940 596312 173164 596340
rect 126940 596300 126946 596312
rect 173158 596300 173164 596312
rect 173216 596300 173222 596352
rect 188614 596300 188620 596352
rect 188672 596340 188678 596352
rect 202874 596340 202880 596352
rect 188672 596312 202880 596340
rect 188672 596300 188678 596312
rect 202874 596300 202880 596312
rect 202932 596300 202938 596352
rect 211062 596300 211068 596352
rect 211120 596340 211126 596352
rect 283098 596340 283104 596352
rect 211120 596312 283104 596340
rect 211120 596300 211126 596312
rect 283098 596300 283104 596312
rect 283156 596300 283162 596352
rect 284478 596300 284484 596352
rect 284536 596340 284542 596352
rect 322934 596340 322940 596352
rect 284536 596312 322940 596340
rect 284536 596300 284542 596312
rect 322934 596300 322940 596312
rect 322992 596300 322998 596352
rect 406470 596300 406476 596352
rect 406528 596340 406534 596352
rect 434714 596340 434720 596352
rect 406528 596312 434720 596340
rect 406528 596300 406534 596312
rect 434714 596300 434720 596312
rect 434772 596300 434778 596352
rect 79778 596232 79784 596284
rect 79836 596272 79842 596284
rect 94038 596272 94044 596284
rect 79836 596244 94044 596272
rect 79836 596232 79842 596244
rect 94038 596232 94044 596244
rect 94096 596232 94102 596284
rect 121362 596232 121368 596284
rect 121420 596272 121426 596284
rect 171962 596272 171968 596284
rect 121420 596244 171968 596272
rect 121420 596232 121426 596244
rect 171962 596232 171968 596244
rect 172020 596232 172026 596284
rect 188706 596232 188712 596284
rect 188764 596272 188770 596284
rect 204346 596272 204352 596284
rect 188764 596244 204352 596272
rect 188764 596232 188770 596244
rect 204346 596232 204352 596244
rect 204404 596232 204410 596284
rect 284386 596232 284392 596284
rect 284444 596272 284450 596284
rect 324406 596272 324412 596284
rect 284444 596244 324412 596272
rect 284444 596232 284450 596244
rect 324406 596232 324412 596244
rect 324464 596232 324470 596284
rect 409322 596232 409328 596284
rect 409380 596272 409386 596284
rect 444374 596272 444380 596284
rect 409380 596244 444380 596272
rect 409380 596232 409386 596244
rect 444374 596232 444380 596244
rect 444432 596232 444438 596284
rect 79962 596164 79968 596216
rect 80020 596204 80026 596216
rect 95234 596204 95240 596216
rect 80020 596176 95240 596204
rect 80020 596164 80026 596176
rect 95234 596164 95240 596176
rect 95292 596164 95298 596216
rect 115842 596164 115848 596216
rect 115900 596204 115906 596216
rect 172146 596204 172152 596216
rect 115900 596176 172152 596204
rect 115900 596164 115906 596176
rect 172146 596164 172152 596176
rect 172204 596164 172210 596216
rect 188522 596164 188528 596216
rect 188580 596204 188586 596216
rect 204254 596204 204260 596216
rect 188580 596176 204260 596204
rect 188580 596164 188586 596176
rect 204254 596164 204260 596176
rect 204312 596164 204318 596216
rect 207106 596164 207112 596216
rect 207164 596204 207170 596216
rect 280982 596204 280988 596216
rect 207164 596176 280988 596204
rect 207164 596164 207170 596176
rect 280982 596164 280988 596176
rect 281040 596164 281046 596216
rect 299382 596164 299388 596216
rect 299440 596204 299446 596216
rect 311894 596204 311900 596216
rect 299440 596176 311900 596204
rect 299440 596164 299446 596176
rect 311894 596164 311900 596176
rect 311952 596164 311958 596216
rect 409230 596164 409236 596216
rect 409288 596204 409294 596216
rect 455414 596204 455420 596216
rect 409288 596176 455420 596204
rect 409288 596164 409294 596176
rect 455414 596164 455420 596176
rect 455472 596164 455478 596216
rect 282178 592628 282184 592680
rect 282236 592668 282242 592680
rect 440234 592668 440240 592680
rect 282236 592640 440240 592668
rect 282236 592628 282242 592640
rect 440234 592628 440240 592640
rect 440292 592628 440298 592680
rect 284938 590656 284944 590708
rect 284996 590696 285002 590708
rect 580166 590696 580172 590708
rect 284996 590668 580172 590696
rect 284996 590656 285002 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 289078 589908 289084 589960
rect 289136 589948 289142 589960
rect 329834 589948 329840 589960
rect 289136 589920 329840 589948
rect 289136 589908 289142 589920
rect 329834 589908 329840 589920
rect 329892 589908 329898 589960
rect 287698 588616 287704 588668
rect 287756 588656 287762 588668
rect 324314 588656 324320 588668
rect 287756 588628 324320 588656
rect 287756 588616 287762 588628
rect 324314 588616 324320 588628
rect 324372 588616 324378 588668
rect 282270 588548 282276 588600
rect 282328 588588 282334 588600
rect 449894 588588 449900 588600
rect 282328 588560 449900 588588
rect 282328 588548 282334 588560
rect 449894 588548 449900 588560
rect 449952 588548 449958 588600
rect 78306 587120 78312 587172
rect 78364 587160 78370 587172
rect 186774 587160 186780 587172
rect 78364 587132 186780 587160
rect 78364 587120 78370 587132
rect 186774 587120 186780 587132
rect 186832 587120 186838 587172
rect 286410 587120 286416 587172
rect 286468 587160 286474 587172
rect 360194 587160 360200 587172
rect 286468 587132 360200 587160
rect 286468 587120 286474 587132
rect 360194 587120 360200 587132
rect 360252 587120 360258 587172
rect 298830 585828 298836 585880
rect 298888 585868 298894 585880
rect 354674 585868 354680 585880
rect 298888 585840 354680 585868
rect 298888 585828 298894 585840
rect 354674 585828 354680 585840
rect 354732 585828 354738 585880
rect 298002 585760 298008 585812
rect 298060 585800 298066 585812
rect 407666 585800 407672 585812
rect 298060 585772 407672 585800
rect 298060 585760 298066 585772
rect 407666 585760 407672 585772
rect 407724 585760 407730 585812
rect 297174 585148 297180 585200
rect 297232 585188 297238 585200
rect 298002 585188 298008 585200
rect 297232 585160 298008 585188
rect 297232 585148 297238 585160
rect 298002 585148 298008 585160
rect 298060 585148 298066 585200
rect 293310 584400 293316 584452
rect 293368 584440 293374 584452
rect 349154 584440 349160 584452
rect 293368 584412 349160 584440
rect 293368 584400 293374 584412
rect 349154 584400 349160 584412
rect 349212 584400 349218 584452
rect 283558 582972 283564 583024
rect 283616 583012 283622 583024
rect 339494 583012 339500 583024
rect 283616 582984 339500 583012
rect 283616 582972 283622 582984
rect 339494 582972 339500 582984
rect 339552 582972 339558 583024
rect 226242 581612 226248 581664
rect 226300 581652 226306 581664
rect 281718 581652 281724 581664
rect 226300 581624 281724 581652
rect 226300 581612 226306 581624
rect 281718 581612 281724 581624
rect 281776 581612 281782 581664
rect 289170 581612 289176 581664
rect 289228 581652 289234 581664
rect 345014 581652 345020 581664
rect 289228 581624 345020 581652
rect 289228 581612 289234 581624
rect 345014 581612 345020 581624
rect 345072 581612 345078 581664
rect 251082 580524 251088 580576
rect 251140 580564 251146 580576
rect 282086 580564 282092 580576
rect 251140 580536 282092 580564
rect 251140 580524 251146 580536
rect 282086 580524 282092 580536
rect 282144 580524 282150 580576
rect 245562 580456 245568 580508
rect 245620 580496 245626 580508
rect 281074 580496 281080 580508
rect 245620 580468 281080 580496
rect 245620 580456 245626 580468
rect 281074 580456 281080 580468
rect 281132 580456 281138 580508
rect 241422 580388 241428 580440
rect 241480 580428 241486 580440
rect 281810 580428 281816 580440
rect 241480 580400 281816 580428
rect 241480 580388 241486 580400
rect 281810 580388 281816 580400
rect 281868 580388 281874 580440
rect 189994 580320 190000 580372
rect 190052 580360 190058 580372
rect 215294 580360 215300 580372
rect 190052 580332 215300 580360
rect 190052 580320 190058 580332
rect 215294 580320 215300 580332
rect 215352 580320 215358 580372
rect 235902 580320 235908 580372
rect 235960 580360 235966 580372
rect 281902 580360 281908 580372
rect 235960 580332 281908 580360
rect 235960 580320 235966 580332
rect 281902 580320 281908 580332
rect 281960 580320 281966 580372
rect 285030 580320 285036 580372
rect 285088 580360 285094 580372
rect 335354 580360 335360 580372
rect 285088 580332 335360 580360
rect 285088 580320 285094 580332
rect 335354 580320 335360 580332
rect 335412 580320 335418 580372
rect 106182 580252 106188 580304
rect 106240 580292 106246 580304
rect 172054 580292 172060 580304
rect 106240 580264 172060 580292
rect 106240 580252 106246 580264
rect 172054 580252 172060 580264
rect 172112 580252 172118 580304
rect 189902 580252 189908 580304
rect 189960 580292 189966 580304
rect 219434 580292 219440 580304
rect 189960 580264 219440 580292
rect 189960 580252 189966 580264
rect 219434 580252 219440 580264
rect 219492 580252 219498 580304
rect 231762 580252 231768 580304
rect 231820 580292 231826 580304
rect 281994 580292 282000 580304
rect 231820 580264 282000 580292
rect 231820 580252 231826 580264
rect 281994 580252 282000 580264
rect 282052 580252 282058 580304
rect 282362 580252 282368 580304
rect 282420 580292 282426 580304
rect 459554 580292 459560 580304
rect 282420 580264 459560 580292
rect 282420 580252 282426 580264
rect 459554 580252 459560 580264
rect 459612 580252 459618 580304
rect 516778 576852 516784 576904
rect 516836 576892 516842 576904
rect 580166 576892 580172 576904
rect 516836 576864 580172 576892
rect 516836 576852 516842 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3326 565836 3332 565888
rect 3384 565876 3390 565888
rect 32398 565876 32404 565888
rect 3384 565848 32404 565876
rect 3384 565836 3390 565848
rect 32398 565836 32404 565848
rect 32456 565836 32462 565888
rect 507118 563048 507124 563100
rect 507176 563088 507182 563100
rect 580166 563088 580172 563100
rect 507176 563060 580172 563088
rect 507176 563048 507182 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3142 553392 3148 553444
rect 3200 553432 3206 553444
rect 22738 553432 22744 553444
rect 3200 553404 22744 553432
rect 3200 553392 3206 553404
rect 22738 553392 22744 553404
rect 22796 553392 22802 553444
rect 511258 536800 511264 536852
rect 511316 536840 511322 536852
rect 579890 536840 579896 536852
rect 511316 536812 579896 536840
rect 511316 536800 511322 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 14458 527184 14464 527196
rect 3384 527156 14464 527184
rect 3384 527144 3390 527156
rect 14458 527144 14464 527156
rect 14516 527144 14522 527196
rect 293862 527008 293868 527060
rect 293920 527048 293926 527060
rect 297266 527048 297272 527060
rect 293920 527020 297272 527048
rect 293920 527008 293926 527020
rect 297266 527008 297272 527020
rect 297324 527048 297330 527060
rect 298002 527048 298008 527060
rect 297324 527020 298008 527048
rect 297324 527008 297330 527020
rect 298002 527008 298008 527020
rect 298060 527008 298066 527060
rect 187326 525784 187332 525836
rect 187384 525824 187390 525836
rect 187694 525824 187700 525836
rect 187384 525796 187700 525824
rect 187384 525784 187390 525796
rect 187694 525784 187700 525796
rect 187752 525784 187758 525836
rect 514018 524424 514024 524476
rect 514076 524464 514082 524476
rect 580166 524464 580172 524476
rect 514076 524436 580172 524464
rect 514076 524424 514082 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 502978 510620 502984 510672
rect 503036 510660 503042 510672
rect 580166 510660 580172 510672
rect 503036 510632 580172 510660
rect 503036 510620 503042 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 10318 501004 10324 501016
rect 3292 500976 10324 501004
rect 3292 500964 3298 500976
rect 10318 500964 10324 500976
rect 10376 500964 10382 501016
rect 287790 498788 287796 498840
rect 287848 498828 287854 498840
rect 297082 498828 297088 498840
rect 287848 498800 297088 498828
rect 287848 498788 287854 498800
rect 297082 498788 297088 498800
rect 297140 498788 297146 498840
rect 78490 489812 78496 489864
rect 78548 489852 78554 489864
rect 187694 489852 187700 489864
rect 78548 489824 187700 489852
rect 78548 489812 78554 489824
rect 187694 489812 187700 489824
rect 187752 489812 187758 489864
rect 407758 489852 407764 489864
rect 306346 489824 407764 489852
rect 78306 489744 78312 489796
rect 78364 489784 78370 489796
rect 187510 489784 187516 489796
rect 78364 489756 187516 489784
rect 78364 489744 78370 489756
rect 187510 489744 187516 489756
rect 187568 489744 187574 489796
rect 297634 489744 297640 489796
rect 297692 489784 297698 489796
rect 306346 489784 306374 489824
rect 407758 489812 407764 489824
rect 407816 489812 407822 489864
rect 297692 489756 306374 489784
rect 297692 489744 297698 489756
rect 78122 489676 78128 489728
rect 78180 489716 78186 489728
rect 187142 489716 187148 489728
rect 78180 489688 187148 489716
rect 78180 489676 78186 489688
rect 187142 489676 187148 489688
rect 187200 489676 187206 489728
rect 77754 489608 77760 489660
rect 77812 489648 77818 489660
rect 187326 489648 187332 489660
rect 77812 489620 187332 489648
rect 77812 489608 77818 489620
rect 187326 489608 187332 489620
rect 187384 489608 187390 489660
rect 78030 489540 78036 489592
rect 78088 489580 78094 489592
rect 187050 489580 187056 489592
rect 78088 489552 187056 489580
rect 78088 489540 78094 489552
rect 187050 489540 187056 489552
rect 187108 489540 187114 489592
rect 78398 489472 78404 489524
rect 78456 489512 78462 489524
rect 186958 489512 186964 489524
rect 78456 489484 186964 489512
rect 78456 489472 78462 489484
rect 186958 489472 186964 489484
rect 187016 489472 187022 489524
rect 77846 489404 77852 489456
rect 77904 489444 77910 489456
rect 186866 489444 186872 489456
rect 77904 489416 186872 489444
rect 77904 489404 77910 489416
rect 186866 489404 186872 489416
rect 186924 489404 186930 489456
rect 78582 489336 78588 489388
rect 78640 489376 78646 489388
rect 186774 489376 186780 489388
rect 78640 489348 186780 489376
rect 78640 489336 78646 489348
rect 186774 489336 186780 489348
rect 186832 489336 186838 489388
rect 173342 489200 173348 489252
rect 173400 489240 173406 489252
rect 253566 489240 253572 489252
rect 173400 489212 253572 489240
rect 173400 489200 173406 489212
rect 253566 489200 253572 489212
rect 253624 489200 253630 489252
rect 218054 489132 218060 489184
rect 218112 489172 218118 489184
rect 404998 489172 405004 489184
rect 218112 489144 405004 489172
rect 218112 489132 218118 489144
rect 404998 489132 405004 489144
rect 405056 489132 405062 489184
rect 186866 488656 186872 488708
rect 186924 488696 186930 488708
rect 187602 488696 187608 488708
rect 186924 488668 187608 488696
rect 186924 488656 186930 488668
rect 187602 488656 187608 488668
rect 187660 488656 187666 488708
rect 187050 488588 187056 488640
rect 187108 488628 187114 488640
rect 187418 488628 187424 488640
rect 187108 488600 187424 488628
rect 187108 488588 187114 488600
rect 187418 488588 187424 488600
rect 187476 488588 187482 488640
rect 186958 488520 186964 488572
rect 187016 488560 187022 488572
rect 187234 488560 187240 488572
rect 187016 488532 187240 488560
rect 187016 488520 187022 488532
rect 187234 488520 187240 488532
rect 187292 488520 187298 488572
rect 79870 488452 79876 488504
rect 79928 488492 79934 488504
rect 92934 488492 92940 488504
rect 79928 488464 92940 488492
rect 79928 488452 79934 488464
rect 92934 488452 92940 488464
rect 92992 488492 92998 488504
rect 188614 488492 188620 488504
rect 92992 488464 188620 488492
rect 92992 488452 92998 488464
rect 188614 488452 188620 488464
rect 188672 488452 188678 488504
rect 407942 488452 407948 488504
rect 408000 488492 408006 488504
rect 425054 488492 425060 488504
rect 408000 488464 425060 488492
rect 408000 488452 408006 488464
rect 425054 488452 425060 488464
rect 425112 488452 425118 488504
rect 79778 488384 79784 488436
rect 79836 488424 79842 488436
rect 94222 488424 94228 488436
rect 79836 488396 94228 488424
rect 79836 488384 79842 488396
rect 94222 488384 94228 488396
rect 94280 488424 94286 488436
rect 188522 488424 188528 488436
rect 94280 488396 188528 488424
rect 94280 488384 94286 488396
rect 188522 488384 188528 488396
rect 188580 488424 188586 488436
rect 204438 488424 204444 488436
rect 188580 488396 204444 488424
rect 188580 488384 188586 488396
rect 204438 488384 204444 488396
rect 204496 488384 204502 488436
rect 291930 488384 291936 488436
rect 291988 488424 291994 488436
rect 297818 488424 297824 488436
rect 291988 488396 297824 488424
rect 291988 488384 291994 488396
rect 297818 488384 297824 488396
rect 297876 488424 297882 488436
rect 407850 488424 407856 488436
rect 297876 488396 407856 488424
rect 297876 488384 297882 488396
rect 407850 488384 407856 488396
rect 407908 488384 407914 488436
rect 408034 488384 408040 488436
rect 408092 488424 408098 488436
rect 423674 488424 423680 488436
rect 408092 488396 423680 488424
rect 408092 488384 408098 488396
rect 423674 488384 423680 488396
rect 423732 488384 423738 488436
rect 79962 488316 79968 488368
rect 80020 488356 80026 488368
rect 95326 488356 95332 488368
rect 80020 488328 95332 488356
rect 80020 488316 80026 488328
rect 95326 488316 95332 488328
rect 95384 488356 95390 488368
rect 95384 488328 180794 488356
rect 95384 488316 95390 488328
rect 180766 488152 180794 488328
rect 297266 488316 297272 488368
rect 297324 488356 297330 488368
rect 407482 488356 407488 488368
rect 297324 488328 407488 488356
rect 297324 488316 297330 488328
rect 407482 488316 407488 488328
rect 407540 488316 407546 488368
rect 408126 488316 408132 488368
rect 408184 488356 408190 488368
rect 422570 488356 422576 488368
rect 408184 488328 422576 488356
rect 408184 488316 408190 488328
rect 422570 488316 422576 488328
rect 422628 488316 422634 488368
rect 299198 488248 299204 488300
rect 299256 488288 299262 488300
rect 314286 488288 314292 488300
rect 299256 488260 314292 488288
rect 299256 488248 299262 488260
rect 314286 488248 314292 488260
rect 314344 488288 314350 488300
rect 408034 488288 408040 488300
rect 314344 488260 408040 488288
rect 314344 488248 314350 488260
rect 408034 488248 408040 488260
rect 408092 488248 408098 488300
rect 188614 488180 188620 488232
rect 188672 488220 188678 488232
rect 202874 488220 202880 488232
rect 188672 488192 202880 488220
rect 188672 488180 188678 488192
rect 202874 488180 202880 488192
rect 202932 488180 202938 488232
rect 299290 488180 299296 488232
rect 299348 488220 299354 488232
rect 315390 488220 315396 488232
rect 299348 488192 315396 488220
rect 299348 488180 299354 488192
rect 315390 488180 315396 488192
rect 315448 488220 315454 488232
rect 407942 488220 407948 488232
rect 315448 488192 407948 488220
rect 315448 488180 315454 488192
rect 407942 488180 407948 488192
rect 408000 488180 408006 488232
rect 188706 488152 188712 488164
rect 180766 488124 188712 488152
rect 188706 488112 188712 488124
rect 188764 488152 188770 488164
rect 204898 488152 204904 488164
rect 188764 488124 204904 488152
rect 188764 488112 188770 488124
rect 204898 488112 204904 488124
rect 204956 488112 204962 488164
rect 297910 488112 297916 488164
rect 297968 488152 297974 488164
rect 408310 488152 408316 488164
rect 297968 488124 408316 488152
rect 297968 488112 297974 488124
rect 408310 488112 408316 488124
rect 408368 488112 408374 488164
rect 188798 488044 188804 488096
rect 188856 488084 188862 488096
rect 220078 488084 220084 488096
rect 188856 488056 220084 488084
rect 188856 488044 188862 488056
rect 220078 488044 220084 488056
rect 220136 488044 220142 488096
rect 104802 487976 104808 488028
rect 104860 488016 104866 488028
rect 214834 488016 214840 488028
rect 104860 487988 214840 488016
rect 104860 487976 104866 487988
rect 214834 487976 214840 487988
rect 214892 487976 214898 488028
rect 230566 487976 230572 488028
rect 230624 488016 230630 488028
rect 287790 488016 287796 488028
rect 230624 487988 287796 488016
rect 230624 487976 230630 487988
rect 287790 487976 287796 487988
rect 287848 487976 287854 488028
rect 103422 487908 103428 487960
rect 103480 487948 103486 487960
rect 213730 487948 213736 487960
rect 103480 487920 213736 487948
rect 103480 487908 103486 487920
rect 213730 487908 213736 487920
rect 213788 487908 213794 487960
rect 219802 487908 219808 487960
rect 219860 487948 219866 487960
rect 281534 487948 281540 487960
rect 219860 487920 281540 487948
rect 219860 487908 219866 487920
rect 281534 487908 281540 487920
rect 281592 487908 281598 487960
rect 105722 487840 105728 487892
rect 105780 487880 105786 487892
rect 215386 487880 215392 487892
rect 105780 487852 215392 487880
rect 105780 487840 105786 487852
rect 215386 487840 215392 487852
rect 215444 487840 215450 487892
rect 232498 487840 232504 487892
rect 232556 487880 232562 487892
rect 299198 487880 299204 487892
rect 232556 487852 299204 487880
rect 232556 487840 232562 487852
rect 299198 487840 299204 487852
rect 299256 487840 299262 487892
rect 101122 487772 101128 487824
rect 101180 487812 101186 487824
rect 211154 487812 211160 487824
rect 101180 487784 211160 487812
rect 101180 487772 101186 487784
rect 211154 487772 211160 487784
rect 211212 487812 211218 487824
rect 212442 487812 212448 487824
rect 211212 487784 212448 487812
rect 211212 487772 211218 487784
rect 212442 487772 212448 487784
rect 212500 487772 212506 487824
rect 232590 487772 232596 487824
rect 232648 487812 232654 487824
rect 299290 487812 299296 487824
rect 232648 487784 299296 487812
rect 232648 487772 232654 487784
rect 299290 487772 299296 487784
rect 299348 487772 299354 487824
rect 312538 487772 312544 487824
rect 312596 487812 312602 487824
rect 312998 487812 313004 487824
rect 312596 487784 313004 487812
rect 312596 487772 312602 487784
rect 312998 487772 313004 487784
rect 313056 487812 313062 487824
rect 408126 487812 408132 487824
rect 313056 487784 408132 487812
rect 313056 487772 313062 487784
rect 408126 487772 408132 487784
rect 408184 487772 408190 487824
rect 319622 487636 319628 487688
rect 319680 487676 319686 487688
rect 427814 487676 427820 487688
rect 319680 487648 427820 487676
rect 319680 487636 319686 487648
rect 427814 487636 427820 487648
rect 427872 487636 427878 487688
rect 326338 487568 326344 487620
rect 326396 487608 326402 487620
rect 434714 487608 434720 487620
rect 326396 487580 434720 487608
rect 326396 487568 326402 487580
rect 434714 487568 434720 487580
rect 434772 487568 434778 487620
rect 318058 487500 318064 487552
rect 318116 487540 318122 487552
rect 426434 487540 426440 487552
rect 318116 487512 426440 487540
rect 318116 487500 318122 487512
rect 426434 487500 426440 487512
rect 426492 487500 426498 487552
rect 204438 487432 204444 487484
rect 204496 487472 204502 487484
rect 222838 487472 222844 487484
rect 204496 487444 222844 487472
rect 204496 487432 204502 487444
rect 222838 487432 222844 487444
rect 222896 487432 222902 487484
rect 322934 487432 322940 487484
rect 322992 487472 322998 487484
rect 433334 487472 433340 487484
rect 322992 487444 433340 487472
rect 322992 487432 322998 487444
rect 433334 487432 433340 487444
rect 433392 487432 433398 487484
rect 102410 487364 102416 487416
rect 102468 487404 102474 487416
rect 211798 487404 211804 487416
rect 102468 487376 211804 487404
rect 102468 487364 102474 487376
rect 211798 487364 211804 487376
rect 211856 487364 211862 487416
rect 212442 487364 212448 487416
rect 212500 487404 212506 487416
rect 226978 487404 226984 487416
rect 212500 487376 226984 487404
rect 212500 487364 212506 487376
rect 226978 487364 226984 487376
rect 227036 487364 227042 487416
rect 324958 487364 324964 487416
rect 325016 487404 325022 487416
rect 434714 487404 434720 487416
rect 325016 487376 434720 487404
rect 325016 487364 325022 487376
rect 434714 487364 434720 487376
rect 434772 487364 434778 487416
rect 100018 487296 100024 487348
rect 100076 487336 100082 487348
rect 210418 487336 210424 487348
rect 100076 487308 210424 487336
rect 100076 487296 100082 487308
rect 210418 487296 210424 487308
rect 210476 487296 210482 487348
rect 214834 487296 214840 487348
rect 214892 487336 214898 487348
rect 229738 487336 229744 487348
rect 214892 487308 229744 487336
rect 214892 487296 214898 487308
rect 229738 487296 229744 487308
rect 229796 487296 229802 487348
rect 320910 487296 320916 487348
rect 320968 487336 320974 487348
rect 430574 487336 430580 487348
rect 320968 487308 430580 487336
rect 320968 487296 320974 487308
rect 430574 487296 430580 487308
rect 430632 487296 430638 487348
rect 98914 487228 98920 487280
rect 98972 487268 98978 487280
rect 209038 487268 209044 487280
rect 98972 487240 209044 487268
rect 98972 487228 98978 487240
rect 209038 487228 209044 487240
rect 209096 487228 209102 487280
rect 213730 487228 213736 487280
rect 213788 487268 213794 487280
rect 229830 487268 229836 487280
rect 213788 487240 229836 487268
rect 213788 487228 213794 487240
rect 229830 487228 229836 487240
rect 229888 487228 229894 487280
rect 320082 487228 320088 487280
rect 320140 487268 320146 487280
rect 429194 487268 429200 487280
rect 320140 487240 429200 487268
rect 320140 487228 320146 487240
rect 429194 487228 429200 487240
rect 429252 487228 429258 487280
rect 97810 487160 97816 487212
rect 97868 487200 97874 487212
rect 207658 487200 207664 487212
rect 97868 487172 207664 487200
rect 97868 487160 97874 487172
rect 207658 487160 207664 487172
rect 207716 487160 207722 487212
rect 215386 487160 215392 487212
rect 215444 487200 215450 487212
rect 244918 487200 244924 487212
rect 215444 487172 244924 487200
rect 215444 487160 215450 487172
rect 244918 487160 244924 487172
rect 244976 487160 244982 487212
rect 321554 487160 321560 487212
rect 321612 487200 321618 487212
rect 322198 487200 322204 487212
rect 321612 487172 322204 487200
rect 321612 487160 321618 487172
rect 322198 487160 322204 487172
rect 322256 487200 322262 487212
rect 432138 487200 432144 487212
rect 322256 487172 432144 487200
rect 322256 487160 322262 487172
rect 432138 487160 432144 487172
rect 432196 487160 432202 487212
rect 457438 487160 457444 487212
rect 457496 487200 457502 487212
rect 465074 487200 465080 487212
rect 457496 487172 465080 487200
rect 457496 487160 457502 487172
rect 465074 487160 465080 487172
rect 465132 487160 465138 487212
rect 299382 487092 299388 487144
rect 299440 487132 299446 487144
rect 311894 487132 311900 487144
rect 299440 487104 311900 487132
rect 299440 487092 299446 487104
rect 311894 487092 311900 487104
rect 311952 487132 311958 487144
rect 312538 487132 312544 487144
rect 311952 487104 312544 487132
rect 311952 487092 311958 487104
rect 312538 487092 312544 487104
rect 312596 487092 312602 487144
rect 243538 486616 243544 486668
rect 243596 486656 243602 486668
rect 322934 486656 322940 486668
rect 243596 486628 322940 486656
rect 243596 486616 243602 486628
rect 322934 486616 322940 486628
rect 322992 486616 322998 486668
rect 172238 486548 172244 486600
rect 172296 486588 172302 486600
rect 254854 486588 254860 486600
rect 172296 486560 254860 486588
rect 172296 486548 172302 486560
rect 254854 486548 254860 486560
rect 254912 486548 254918 486600
rect 187694 486480 187700 486532
rect 187752 486520 187758 486532
rect 235258 486520 235264 486532
rect 187752 486492 235264 486520
rect 187752 486480 187758 486492
rect 235258 486480 235264 486492
rect 235316 486480 235322 486532
rect 253934 486480 253940 486532
rect 253992 486520 253998 486532
rect 409414 486520 409420 486532
rect 253992 486492 409420 486520
rect 253992 486480 253998 486492
rect 409414 486480 409420 486492
rect 409472 486480 409478 486532
rect 216766 486412 216772 486464
rect 216824 486452 216830 486464
rect 542354 486452 542360 486464
rect 216824 486424 542360 486452
rect 216824 486412 216830 486424
rect 542354 486412 542360 486424
rect 542412 486412 542418 486464
rect 297266 486004 297272 486056
rect 297324 486044 297330 486056
rect 297726 486044 297732 486056
rect 297324 486016 297732 486044
rect 297324 486004 297330 486016
rect 297726 486004 297732 486016
rect 297784 486004 297790 486056
rect 296806 485936 296812 485988
rect 296864 485976 296870 485988
rect 297910 485976 297916 485988
rect 296864 485948 297916 485976
rect 296864 485936 296870 485948
rect 297910 485936 297916 485948
rect 297968 485936 297974 485988
rect 243630 485800 243636 485852
rect 243688 485840 243694 485852
rect 244642 485840 244648 485852
rect 243688 485812 244648 485840
rect 243688 485800 243694 485812
rect 244642 485800 244648 485812
rect 244700 485800 244706 485852
rect 240778 485120 240784 485172
rect 240836 485160 240842 485172
rect 320910 485160 320916 485172
rect 240836 485132 320916 485160
rect 240836 485120 240842 485132
rect 320910 485120 320916 485132
rect 320968 485120 320974 485172
rect 173250 485052 173256 485104
rect 173308 485092 173314 485104
rect 247218 485092 247224 485104
rect 173308 485064 247224 485092
rect 173308 485052 173314 485064
rect 247218 485052 247224 485064
rect 247276 485052 247282 485104
rect 248414 485052 248420 485104
rect 248472 485092 248478 485104
rect 409322 485092 409328 485104
rect 248472 485064 409328 485092
rect 248472 485052 248478 485064
rect 409322 485052 409328 485064
rect 409380 485052 409386 485104
rect 221458 484372 221464 484424
rect 221516 484412 221522 484424
rect 580166 484412 580172 484424
rect 221516 484384 580172 484412
rect 221516 484372 221522 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 251634 483692 251640 483744
rect 251692 483732 251698 483744
rect 409230 483732 409236 483744
rect 251692 483704 409236 483732
rect 251692 483692 251698 483704
rect 409230 483692 409236 483704
rect 409288 483692 409294 483744
rect 216950 483624 216956 483676
rect 217008 483664 217014 483676
rect 580258 483664 580264 483676
rect 217008 483636 580264 483664
rect 217008 483624 217014 483636
rect 580258 483624 580264 483636
rect 580316 483624 580322 483676
rect 242158 482400 242164 482452
rect 242216 482440 242222 482452
rect 321554 482440 321560 482452
rect 242216 482412 321560 482440
rect 242216 482400 242222 482412
rect 321554 482400 321560 482412
rect 321612 482400 321618 482452
rect 105998 482332 106004 482384
rect 106056 482372 106062 482384
rect 234614 482372 234620 482384
rect 106056 482344 234620 482372
rect 106056 482332 106062 482344
rect 234614 482332 234620 482344
rect 234672 482332 234678 482384
rect 246390 482332 246396 482384
rect 246448 482372 246454 482384
rect 360194 482372 360200 482384
rect 246448 482344 360200 482372
rect 246448 482332 246454 482344
rect 360194 482332 360200 482344
rect 360252 482332 360258 482384
rect 216674 482264 216680 482316
rect 216732 482304 216738 482316
rect 501598 482304 501604 482316
rect 216732 482276 501604 482304
rect 216732 482264 216738 482276
rect 501598 482264 501604 482276
rect 501656 482264 501662 482316
rect 173158 481040 173164 481092
rect 173216 481080 173222 481092
rect 250990 481080 250996 481092
rect 173216 481052 250996 481080
rect 173216 481040 173222 481052
rect 250990 481040 250996 481052
rect 251048 481040 251054 481092
rect 236086 480972 236092 481024
rect 236144 481012 236150 481024
rect 434714 481012 434720 481024
rect 236144 480984 434720 481012
rect 236144 480972 236150 480984
rect 434714 480972 434720 480984
rect 434772 480972 434778 481024
rect 215294 480904 215300 480956
rect 215352 480944 215358 480956
rect 516778 480944 516784 480956
rect 215352 480916 516784 480944
rect 215352 480904 215358 480916
rect 516778 480904 516784 480916
rect 516836 480904 516842 480956
rect 238110 479680 238116 479732
rect 238168 479720 238174 479732
rect 319622 479720 319628 479732
rect 238168 479692 319628 479720
rect 238168 479680 238174 479692
rect 319622 479680 319628 479692
rect 319680 479680 319686 479732
rect 238846 479612 238852 479664
rect 238904 479652 238910 479664
rect 339494 479652 339500 479664
rect 238904 479624 339500 479652
rect 238904 479612 238910 479624
rect 339494 479612 339500 479624
rect 339552 479612 339558 479664
rect 126882 479544 126888 479596
rect 126940 479584 126946 479596
rect 240870 479584 240876 479596
rect 126940 479556 240876 479584
rect 126940 479544 126946 479556
rect 240870 479544 240876 479556
rect 240928 479544 240934 479596
rect 215478 479476 215484 479528
rect 215536 479516 215542 479528
rect 514018 479516 514024 479528
rect 215536 479488 514024 479516
rect 215536 479476 215542 479488
rect 514018 479476 514024 479488
rect 514076 479476 514082 479528
rect 172146 478320 172152 478372
rect 172204 478360 172210 478372
rect 248506 478360 248512 478372
rect 172204 478332 248512 478360
rect 172204 478320 172210 478332
rect 248506 478320 248512 478332
rect 248564 478320 248570 478372
rect 246482 478252 246488 478304
rect 246540 478292 246546 478304
rect 354674 478292 354680 478304
rect 246540 478264 354680 478292
rect 246540 478252 246546 478264
rect 354674 478252 354680 478264
rect 354732 478252 354738 478304
rect 246758 478184 246764 478236
rect 246816 478224 246822 478236
rect 406470 478224 406476 478236
rect 246816 478196 406476 478224
rect 246816 478184 246822 478196
rect 406470 478184 406476 478196
rect 406528 478184 406534 478236
rect 218238 478116 218244 478168
rect 218296 478156 218302 478168
rect 395338 478156 395344 478168
rect 218296 478128 395344 478156
rect 218296 478116 218302 478128
rect 395338 478116 395344 478128
rect 395396 478116 395402 478168
rect 293402 477476 293408 477488
rect 238726 477448 293408 477476
rect 235258 477368 235264 477420
rect 235316 477408 235322 477420
rect 238726 477408 238754 477448
rect 293402 477436 293408 477448
rect 293460 477436 293466 477488
rect 235316 477380 238754 477408
rect 235316 477368 235322 477380
rect 218146 476824 218152 476876
rect 218204 476864 218210 476876
rect 403618 476864 403624 476876
rect 218204 476836 403624 476864
rect 218204 476824 218210 476836
rect 403618 476824 403624 476836
rect 403676 476824 403682 476876
rect 210418 476756 210424 476808
rect 210476 476796 210482 476808
rect 239398 476796 239404 476808
rect 210476 476768 239404 476796
rect 210476 476756 210482 476768
rect 239398 476756 239404 476768
rect 239456 476756 239462 476808
rect 241606 476756 241612 476808
rect 241664 476796 241670 476808
rect 459554 476796 459560 476808
rect 241664 476768 459560 476796
rect 241664 476756 241670 476768
rect 459554 476756 459560 476768
rect 459612 476756 459618 476808
rect 234798 476076 234804 476128
rect 234856 476116 234862 476128
rect 235258 476116 235264 476128
rect 234856 476088 235264 476116
rect 234856 476076 234862 476088
rect 235258 476076 235264 476088
rect 235316 476076 235322 476128
rect 244366 476008 244372 476060
rect 244424 476048 244430 476060
rect 244918 476048 244924 476060
rect 244424 476020 244924 476048
rect 244424 476008 244430 476020
rect 244918 476008 244924 476020
rect 244976 476048 244982 476060
rect 326338 476048 326344 476060
rect 244976 476020 326344 476048
rect 244976 476008 244982 476020
rect 326338 476008 326344 476020
rect 326396 476008 326402 476060
rect 236270 475396 236276 475448
rect 236328 475436 236334 475448
rect 329834 475436 329840 475448
rect 236328 475408 329840 475436
rect 236328 475396 236334 475408
rect 329834 475396 329840 475408
rect 329892 475396 329898 475448
rect 217134 475328 217140 475380
rect 217192 475368 217198 475380
rect 527174 475368 527180 475380
rect 217192 475340 527180 475368
rect 217192 475328 217198 475340
rect 527174 475328 527180 475340
rect 527232 475328 527238 475380
rect 3234 474716 3240 474768
rect 3292 474756 3298 474768
rect 40678 474756 40684 474768
rect 3292 474728 40684 474756
rect 3292 474716 3298 474728
rect 40678 474716 40684 474728
rect 40736 474716 40742 474768
rect 235902 474648 235908 474700
rect 235960 474688 235966 474700
rect 240962 474688 240968 474700
rect 235960 474660 240968 474688
rect 235960 474648 235966 474660
rect 240962 474648 240968 474660
rect 241020 474648 241026 474700
rect 241422 474648 241428 474700
rect 241480 474688 241486 474700
rect 242250 474688 242256 474700
rect 241480 474660 242256 474688
rect 241480 474648 241486 474660
rect 242250 474648 242256 474660
rect 242308 474648 242314 474700
rect 244918 474104 244924 474156
rect 244976 474144 244982 474156
rect 324958 474144 324964 474156
rect 244976 474116 324964 474144
rect 244976 474104 244982 474116
rect 324958 474104 324964 474116
rect 325016 474104 325022 474156
rect 77938 474036 77944 474088
rect 77996 474076 78002 474088
rect 229922 474076 229928 474088
rect 77996 474048 229928 474076
rect 77996 474036 78002 474048
rect 229922 474036 229928 474048
rect 229980 474036 229986 474088
rect 237926 474036 237932 474088
rect 237984 474076 237990 474088
rect 335354 474076 335360 474088
rect 237984 474048 335360 474076
rect 237984 474036 237990 474048
rect 335354 474036 335360 474048
rect 335412 474036 335418 474088
rect 215662 473968 215668 474020
rect 215720 474008 215726 474020
rect 512638 474008 512644 474020
rect 215720 473980 512644 474008
rect 215720 473968 215726 473980
rect 512638 473968 512644 473980
rect 512696 473968 512702 474020
rect 216582 472744 216588 472796
rect 216640 472784 216646 472796
rect 235534 472784 235540 472796
rect 216640 472756 235540 472784
rect 216640 472744 216646 472756
rect 235534 472744 235540 472756
rect 235592 472744 235598 472796
rect 236638 472744 236644 472796
rect 236696 472784 236702 472796
rect 318058 472784 318064 472796
rect 236696 472756 318064 472784
rect 236696 472744 236702 472756
rect 318058 472744 318064 472756
rect 318116 472744 318122 472796
rect 32398 472676 32404 472728
rect 32456 472716 32462 472728
rect 224310 472716 224316 472728
rect 32456 472688 224316 472716
rect 32456 472676 32462 472688
rect 224310 472676 224316 472688
rect 224368 472676 224374 472728
rect 238018 472676 238024 472728
rect 238076 472716 238082 472728
rect 324314 472716 324320 472728
rect 238076 472688 324320 472716
rect 238076 472676 238082 472688
rect 324314 472676 324320 472688
rect 324372 472676 324378 472728
rect 215386 472608 215392 472660
rect 215444 472648 215450 472660
rect 511258 472648 511264 472660
rect 215444 472620 511264 472648
rect 215444 472608 215450 472620
rect 511258 472608 511264 472620
rect 511316 472608 511322 472660
rect 211798 471928 211804 471980
rect 211856 471968 211862 471980
rect 241698 471968 241704 471980
rect 211856 471940 241704 471968
rect 211856 471928 211862 471940
rect 241698 471928 241704 471940
rect 241756 471968 241762 471980
rect 242158 471968 242164 471980
rect 241756 471940 242164 471968
rect 241756 471928 241762 471940
rect 242158 471928 242164 471940
rect 242216 471928 242222 471980
rect 40678 471248 40684 471300
rect 40736 471288 40742 471300
rect 224494 471288 224500 471300
rect 40736 471260 224500 471288
rect 40736 471248 40742 471260
rect 224494 471248 224500 471260
rect 224552 471248 224558 471300
rect 237466 471248 237472 471300
rect 237524 471288 237530 471300
rect 440234 471288 440240 471300
rect 237524 471260 440240 471288
rect 237524 471248 237530 471260
rect 440234 471248 440240 471260
rect 440292 471248 440298 471300
rect 214006 470568 214012 470620
rect 214064 470608 214070 470620
rect 579982 470608 579988 470620
rect 214064 470580 579988 470608
rect 214064 470568 214070 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 207658 470500 207664 470552
rect 207716 470540 207722 470552
rect 236638 470540 236644 470552
rect 207716 470512 236644 470540
rect 207716 470500 207722 470512
rect 236638 470500 236644 470512
rect 236696 470500 236702 470552
rect 10318 469888 10324 469940
rect 10376 469928 10382 469940
rect 224678 469928 224684 469940
rect 10376 469900 224684 469928
rect 10376 469888 10382 469900
rect 224678 469888 224684 469900
rect 224736 469888 224742 469940
rect 239030 469888 239036 469940
rect 239088 469928 239094 469940
rect 449894 469928 449900 469940
rect 239088 469900 449900 469928
rect 239088 469888 239094 469900
rect 449894 469888 449900 469900
rect 449952 469888 449958 469940
rect 217318 469820 217324 469872
rect 217376 469860 217382 469872
rect 509878 469860 509884 469872
rect 217376 469832 509884 469860
rect 217376 469820 217382 469832
rect 509878 469820 509884 469832
rect 509936 469820 509942 469872
rect 219618 468596 219624 468648
rect 219676 468636 219682 468648
rect 296070 468636 296076 468648
rect 219676 468608 296076 468636
rect 219676 468596 219682 468608
rect 296070 468596 296076 468608
rect 296128 468596 296134 468648
rect 218330 468528 218336 468580
rect 218388 468568 218394 468580
rect 399478 468568 399484 468580
rect 218388 468540 399484 468568
rect 218388 468528 218394 468540
rect 399478 468528 399484 468540
rect 399536 468528 399542 468580
rect 22738 468460 22744 468512
rect 22796 468500 22802 468512
rect 223758 468500 223764 468512
rect 22796 468472 223764 468500
rect 22796 468460 22802 468472
rect 223758 468460 223764 468472
rect 223816 468460 223822 468512
rect 238754 468460 238760 468512
rect 238812 468500 238818 468512
rect 444374 468500 444380 468512
rect 238812 468472 444380 468500
rect 238812 468460 238818 468472
rect 444374 468460 444380 468472
rect 444432 468460 444438 468512
rect 178678 467236 178684 467288
rect 178736 467276 178742 467288
rect 221366 467276 221372 467288
rect 178736 467248 221372 467276
rect 178736 467236 178742 467248
rect 221366 467236 221372 467248
rect 221424 467236 221430 467288
rect 218422 467168 218428 467220
rect 218480 467208 218486 467220
rect 409138 467208 409144 467220
rect 218480 467180 409144 467208
rect 218480 467168 218486 467180
rect 409138 467168 409144 467180
rect 409196 467168 409202 467220
rect 121362 467100 121368 467152
rect 121420 467140 121426 467152
rect 239490 467140 239496 467152
rect 121420 467112 239496 467140
rect 121420 467100 121426 467112
rect 239490 467100 239496 467112
rect 239548 467100 239554 467152
rect 244550 467100 244556 467152
rect 244608 467140 244614 467152
rect 470594 467140 470600 467152
rect 244608 467112 470600 467140
rect 244608 467100 244614 467112
rect 470594 467100 470600 467112
rect 470652 467100 470658 467152
rect 136542 465808 136548 465860
rect 136600 465848 136606 465860
rect 243354 465848 243360 465860
rect 136600 465820 243360 465848
rect 136600 465808 136606 465820
rect 243354 465808 243360 465820
rect 243412 465808 243418 465860
rect 217502 465740 217508 465792
rect 217560 465780 217566 465792
rect 406378 465780 406384 465792
rect 217560 465752 406384 465780
rect 217560 465740 217566 465752
rect 406378 465740 406384 465752
rect 406436 465740 406442 465792
rect 243078 465672 243084 465724
rect 243136 465712 243142 465724
rect 457438 465712 457444 465724
rect 243136 465684 457444 465712
rect 243136 465672 243142 465684
rect 457438 465672 457444 465684
rect 457496 465672 457502 465724
rect 220722 464516 220728 464568
rect 220780 464556 220786 464568
rect 237006 464556 237012 464568
rect 220780 464528 237012 464556
rect 220780 464516 220786 464528
rect 237006 464516 237012 464528
rect 237064 464516 237070 464568
rect 231486 464448 231492 464500
rect 231544 464488 231550 464500
rect 311894 464488 311900 464500
rect 231544 464460 311900 464488
rect 231544 464448 231550 464460
rect 311894 464448 311900 464460
rect 311952 464448 311958 464500
rect 4062 464380 4068 464432
rect 4120 464420 4126 464432
rect 224218 464420 224224 464432
rect 4120 464392 224224 464420
rect 4120 464380 4126 464392
rect 224218 464380 224224 464392
rect 224276 464380 224282 464432
rect 240318 464380 240324 464432
rect 240376 464420 240382 464432
rect 454678 464420 454684 464432
rect 240376 464392 454684 464420
rect 240376 464380 240382 464392
rect 454678 464380 454684 464392
rect 454736 464380 454742 464432
rect 215846 464312 215852 464364
rect 215904 464352 215910 464364
rect 504358 464352 504364 464364
rect 215904 464324 504364 464352
rect 215904 464312 215910 464324
rect 504358 464312 504364 464324
rect 504416 464312 504422 464364
rect 209038 463632 209044 463684
rect 209096 463672 209102 463684
rect 237558 463672 237564 463684
rect 209096 463644 237564 463672
rect 209096 463632 209102 463644
rect 237558 463632 237564 463644
rect 237616 463672 237622 463684
rect 238110 463672 238116 463684
rect 237616 463644 238116 463672
rect 237616 463632 237622 463644
rect 238110 463632 238116 463644
rect 238168 463632 238174 463684
rect 219710 463156 219716 463208
rect 219768 463196 219774 463208
rect 282914 463196 282920 463208
rect 219768 463168 282920 463196
rect 219768 463156 219774 463168
rect 282914 463156 282920 463168
rect 282972 463156 282978 463208
rect 240502 463088 240508 463140
rect 240560 463128 240566 463140
rect 345014 463128 345020 463140
rect 240560 463100 345020 463128
rect 240560 463088 240566 463100
rect 345014 463088 345020 463100
rect 345072 463088 345078 463140
rect 230750 463020 230756 463072
rect 230808 463060 230814 463072
rect 408218 463060 408224 463072
rect 230808 463032 408224 463060
rect 230808 463020 230814 463032
rect 408218 463020 408224 463032
rect 408276 463020 408282 463072
rect 216858 462952 216864 463004
rect 216916 462992 216922 463004
rect 508498 462992 508504 463004
rect 216916 462964 508504 462992
rect 216916 462952 216922 462964
rect 508498 462952 508504 462964
rect 508556 462952 508562 463004
rect 2866 462340 2872 462392
rect 2924 462380 2930 462392
rect 225598 462380 225604 462392
rect 2924 462352 225604 462380
rect 2924 462340 2930 462352
rect 225598 462340 225604 462352
rect 225656 462340 225662 462392
rect 219894 461796 219900 461848
rect 219952 461836 219958 461848
rect 291838 461836 291844 461848
rect 219952 461808 291844 461836
rect 219952 461796 219958 461808
rect 291838 461796 291844 461808
rect 291896 461796 291902 461848
rect 131022 461728 131028 461780
rect 131080 461768 131086 461780
rect 242066 461768 242072 461780
rect 131080 461740 242072 461768
rect 131080 461728 131086 461740
rect 242066 461728 242072 461740
rect 242124 461728 242130 461780
rect 71774 461660 71780 461712
rect 71832 461700 71838 461712
rect 221550 461700 221556 461712
rect 71832 461672 221556 461700
rect 71832 461660 71838 461672
rect 221550 461660 221556 461672
rect 221608 461660 221614 461712
rect 241790 461660 241796 461712
rect 241848 461700 241854 461712
rect 349154 461700 349160 461712
rect 241848 461672 349160 461700
rect 241848 461660 241854 461672
rect 349154 461660 349160 461672
rect 349212 461660 349218 461712
rect 215754 461592 215760 461644
rect 215812 461632 215818 461644
rect 507118 461632 507124 461644
rect 215812 461604 507124 461632
rect 215812 461592 215818 461604
rect 507118 461592 507124 461604
rect 507176 461592 507182 461644
rect 319438 460884 319444 460896
rect 248386 460856 319444 460884
rect 239398 460776 239404 460828
rect 239456 460816 239462 460828
rect 248386 460816 248414 460856
rect 319438 460844 319444 460856
rect 319496 460844 319502 460896
rect 239456 460788 248414 460816
rect 239456 460776 239462 460788
rect 218606 460300 218612 460352
rect 218664 460340 218670 460352
rect 293218 460340 293224 460352
rect 218664 460312 293224 460340
rect 218664 460300 218670 460312
rect 293218 460300 293224 460312
rect 293276 460300 293282 460352
rect 14458 460232 14464 460284
rect 14516 460272 14522 460284
rect 224034 460272 224040 460284
rect 14516 460244 224040 460272
rect 14516 460232 14522 460244
rect 224034 460232 224040 460244
rect 224092 460232 224098 460284
rect 214190 460164 214196 460216
rect 214248 460204 214254 460216
rect 502978 460204 502984 460216
rect 214248 460176 502984 460204
rect 214248 460164 214254 460176
rect 502978 460164 502984 460176
rect 503036 460164 503042 460216
rect 203518 459484 203524 459536
rect 203576 459524 203582 459536
rect 231578 459524 231584 459536
rect 203576 459496 231584 459524
rect 203576 459484 203582 459496
rect 231578 459484 231584 459496
rect 231636 459484 231642 459536
rect 246298 458940 246304 458992
rect 246356 458980 246362 458992
rect 363138 458980 363144 458992
rect 246356 458952 363144 458980
rect 246356 458940 246362 458952
rect 363138 458940 363144 458952
rect 363196 458940 363202 458992
rect 171962 458872 171968 458924
rect 172020 458912 172026 458924
rect 249794 458912 249800 458924
rect 172020 458884 249800 458912
rect 172020 458872 172026 458884
rect 249794 458872 249800 458884
rect 249852 458872 249858 458924
rect 253290 458872 253296 458924
rect 253348 458912 253354 458924
rect 371510 458912 371516 458924
rect 253348 458884 371516 458912
rect 253348 458872 253354 458884
rect 371510 458872 371516 458884
rect 371568 458872 371574 458924
rect 40034 458804 40040 458856
rect 40092 458844 40098 458856
rect 220998 458844 221004 458856
rect 40092 458816 221004 458844
rect 40092 458804 40098 458816
rect 220998 458804 221004 458816
rect 221056 458804 221062 458856
rect 247034 458804 247040 458856
rect 247092 458844 247098 458856
rect 379882 458844 379888 458856
rect 247092 458816 379888 458844
rect 247092 458804 247098 458816
rect 379882 458804 379888 458816
rect 379940 458804 379946 458856
rect 299382 458736 299388 458788
rect 299440 458776 299446 458788
rect 329650 458776 329656 458788
rect 299440 458748 329656 458776
rect 299440 458736 299446 458748
rect 329650 458736 329656 458748
rect 329708 458736 329714 458788
rect 299474 458668 299480 458720
rect 299532 458708 299538 458720
rect 342530 458708 342536 458720
rect 299532 458680 342536 458708
rect 299532 458668 299538 458680
rect 342530 458668 342536 458680
rect 342588 458668 342594 458720
rect 296070 458600 296076 458652
rect 296128 458640 296134 458652
rect 346394 458640 346400 458652
rect 296128 458612 346400 458640
rect 296128 458600 296134 458612
rect 346394 458600 346400 458612
rect 346452 458600 346458 458652
rect 299566 458532 299572 458584
rect 299624 458572 299630 458584
rect 350902 458572 350908 458584
rect 299624 458544 350908 458572
rect 299624 458532 299630 458544
rect 350902 458532 350908 458544
rect 350960 458532 350966 458584
rect 298738 458464 298744 458516
rect 298796 458504 298802 458516
rect 359274 458504 359280 458516
rect 298796 458476 359280 458504
rect 298796 458464 298802 458476
rect 359274 458464 359280 458476
rect 359332 458464 359338 458516
rect 298002 458396 298008 458448
rect 298060 458436 298066 458448
rect 367646 458436 367652 458448
rect 298060 458408 367652 458436
rect 298060 458396 298066 458408
rect 367646 458396 367652 458408
rect 367704 458396 367710 458448
rect 355778 458328 355784 458380
rect 355836 458368 355842 458380
rect 376018 458368 376024 458380
rect 355836 458340 376024 458368
rect 355836 458328 355842 458340
rect 376018 458328 376024 458340
rect 376076 458328 376082 458380
rect 293218 458260 293224 458312
rect 293276 458300 293282 458312
rect 309042 458300 309048 458312
rect 293276 458272 309048 458300
rect 293276 458260 293282 458272
rect 309042 458260 309048 458272
rect 309100 458260 309106 458312
rect 299658 458192 299664 458244
rect 299716 458232 299722 458244
rect 321278 458232 321284 458244
rect 299716 458204 321284 458232
rect 299716 458192 299722 458204
rect 321278 458192 321284 458204
rect 321336 458192 321342 458244
rect 174538 457512 174544 457564
rect 174596 457552 174602 457564
rect 221274 457552 221280 457564
rect 174596 457524 221280 457552
rect 174596 457512 174602 457524
rect 221274 457512 221280 457524
rect 221332 457512 221338 457564
rect 6914 457444 6920 457496
rect 6972 457484 6978 457496
rect 220814 457484 220820 457496
rect 6972 457456 220820 457484
rect 6972 457444 6978 457456
rect 220814 457444 220820 457456
rect 220872 457444 220878 457496
rect 227346 457444 227352 457496
rect 227404 457484 227410 457496
rect 355778 457484 355784 457496
rect 227404 457456 355784 457484
rect 227404 457444 227410 457456
rect 355778 457444 355784 457456
rect 355836 457444 355842 457496
rect 222930 457240 222936 457292
rect 222988 457280 222994 457292
rect 317414 457280 317420 457292
rect 222988 457252 317420 457280
rect 222988 457240 222994 457252
rect 317414 457240 317420 457252
rect 317472 457240 317478 457292
rect 228450 457172 228456 457224
rect 228508 457212 228514 457224
rect 325786 457212 325792 457224
rect 228508 457184 325792 457212
rect 228508 457172 228514 457184
rect 325786 457172 325792 457184
rect 325844 457172 325850 457224
rect 236362 457104 236368 457156
rect 236420 457144 236426 457156
rect 338022 457144 338028 457156
rect 236420 457116 338028 457144
rect 236420 457104 236426 457116
rect 338022 457104 338028 457116
rect 338080 457104 338086 457156
rect 228358 457036 228364 457088
rect 228416 457076 228422 457088
rect 334158 457076 334164 457088
rect 228416 457048 334164 457076
rect 228416 457036 228422 457048
rect 334158 457036 334164 457048
rect 334216 457036 334222 457088
rect 247126 456968 247132 457020
rect 247184 457008 247190 457020
rect 354766 457008 354772 457020
rect 247184 456980 354772 457008
rect 247184 456968 247190 456980
rect 354766 456968 354772 456980
rect 354824 456968 354830 457020
rect 223022 456900 223028 456952
rect 223080 456940 223086 456952
rect 383746 456940 383752 456952
rect 223080 456912 383752 456940
rect 223080 456900 223086 456912
rect 383746 456900 383752 456912
rect 383804 456900 383810 456952
rect 385494 456872 385500 456884
rect 229066 456844 385500 456872
rect 223850 456764 223856 456816
rect 223908 456804 223914 456816
rect 224310 456804 224316 456816
rect 223908 456776 224316 456804
rect 223908 456764 223914 456776
rect 224310 456764 224316 456776
rect 224368 456804 224374 456816
rect 229066 456804 229094 456844
rect 385494 456832 385500 456844
rect 385552 456832 385558 456884
rect 224368 456776 229094 456804
rect 224368 456764 224374 456776
rect 299014 456764 299020 456816
rect 299072 456804 299078 456816
rect 580166 456804 580172 456816
rect 299072 456776 580172 456804
rect 299072 456764 299078 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 240502 456084 240508 456136
rect 240560 456124 240566 456136
rect 241146 456124 241152 456136
rect 240560 456096 241152 456124
rect 240560 456084 240566 456096
rect 241146 456084 241152 456096
rect 241204 456084 241210 456136
rect 299750 456084 299756 456136
rect 299808 456124 299814 456136
rect 300762 456124 300768 456136
rect 299808 456096 300768 456124
rect 299808 456084 299814 456096
rect 300762 456084 300768 456096
rect 300820 456084 300826 456136
rect 235074 456016 235080 456068
rect 235132 456056 235138 456068
rect 312630 456056 312636 456068
rect 235132 456028 312636 456056
rect 235132 456016 235138 456028
rect 312630 456016 312636 456028
rect 312688 456016 312694 456068
rect 252646 455948 252652 456000
rect 252704 455988 252710 456000
rect 385310 455988 385316 456000
rect 252704 455960 385316 455988
rect 252704 455948 252710 455960
rect 385310 455948 385316 455960
rect 385368 455948 385374 456000
rect 251726 455880 251732 455932
rect 251784 455920 251790 455932
rect 385402 455920 385408 455932
rect 251784 455892 385408 455920
rect 251784 455880 251790 455892
rect 385402 455880 385408 455892
rect 385460 455880 385466 455932
rect 251358 455812 251364 455864
rect 251416 455852 251422 455864
rect 385034 455852 385040 455864
rect 251416 455824 385040 455852
rect 251416 455812 251422 455824
rect 385034 455812 385040 455824
rect 385092 455812 385098 455864
rect 250162 455744 250168 455796
rect 250220 455784 250226 455796
rect 384114 455784 384120 455796
rect 250220 455756 384120 455784
rect 250220 455744 250226 455756
rect 384114 455744 384120 455756
rect 384172 455744 384178 455796
rect 244458 455676 244464 455728
rect 244516 455716 244522 455728
rect 384206 455716 384212 455728
rect 244516 455688 384212 455716
rect 244516 455676 244522 455688
rect 384206 455676 384212 455688
rect 384264 455676 384270 455728
rect 298922 455608 298928 455660
rect 298980 455648 298986 455660
rect 300302 455648 300308 455660
rect 298980 455620 300308 455648
rect 298980 455608 298986 455620
rect 300302 455608 300308 455620
rect 300360 455608 300366 455660
rect 300762 455608 300768 455660
rect 300820 455648 300826 455660
rect 385218 455648 385224 455660
rect 300820 455620 385224 455648
rect 300820 455608 300826 455620
rect 385218 455608 385224 455620
rect 385276 455608 385282 455660
rect 237742 455540 237748 455592
rect 237800 455580 237806 455592
rect 384022 455580 384028 455592
rect 237800 455552 384028 455580
rect 237800 455540 237806 455552
rect 384022 455540 384028 455552
rect 384080 455540 384086 455592
rect 214282 455472 214288 455524
rect 214340 455512 214346 455524
rect 384298 455512 384304 455524
rect 214340 455484 384304 455512
rect 214340 455472 214346 455484
rect 384298 455472 384304 455484
rect 384356 455472 384362 455524
rect 214466 455404 214472 455456
rect 214524 455444 214530 455456
rect 580258 455444 580264 455456
rect 214524 455416 580264 455444
rect 214524 455404 214530 455416
rect 580258 455404 580264 455416
rect 580316 455404 580322 455456
rect 299842 455336 299848 455388
rect 299900 455376 299906 455388
rect 304166 455376 304172 455388
rect 299900 455348 304172 455376
rect 299900 455336 299906 455348
rect 304166 455336 304172 455348
rect 304224 455336 304230 455388
rect 248690 454860 248696 454912
rect 248748 454900 248754 454912
rect 299842 454900 299848 454912
rect 248748 454872 299848 454900
rect 248748 454860 248754 454872
rect 299842 454860 299848 454872
rect 299900 454860 299906 454912
rect 234706 454792 234712 454844
rect 234764 454832 234770 454844
rect 299566 454832 299572 454844
rect 234764 454804 299572 454832
rect 234764 454792 234770 454804
rect 299566 454792 299572 454804
rect 299624 454792 299630 454844
rect 235258 454724 235264 454776
rect 235316 454764 235322 454776
rect 299474 454764 299480 454776
rect 235316 454736 299480 454764
rect 235316 454724 235322 454736
rect 299474 454724 299480 454736
rect 299532 454724 299538 454776
rect 219066 454656 219072 454708
rect 219124 454696 219130 454708
rect 295978 454696 295984 454708
rect 219124 454668 295984 454696
rect 219124 454656 219130 454668
rect 295978 454656 295984 454668
rect 296036 454656 296042 454708
rect 182818 453432 182824 453484
rect 182876 453472 182882 453484
rect 221090 453472 221096 453484
rect 182876 453444 221096 453472
rect 182876 453432 182882 453444
rect 221090 453432 221096 453444
rect 221148 453432 221154 453484
rect 215938 453364 215944 453416
rect 215996 453404 216002 453416
rect 284938 453404 284944 453416
rect 215996 453376 284944 453404
rect 215996 453364 216002 453376
rect 284938 453364 284944 453376
rect 284996 453364 285002 453416
rect 214650 453296 214656 453348
rect 214708 453336 214714 453348
rect 299014 453336 299020 453348
rect 214708 453308 299020 453336
rect 214708 453296 214714 453308
rect 299014 453296 299020 453308
rect 299072 453296 299078 453348
rect 237558 453092 237564 453144
rect 237616 453132 237622 453144
rect 237834 453132 237840 453144
rect 237616 453104 237840 453132
rect 237616 453092 237622 453104
rect 237834 453092 237840 453104
rect 237892 453092 237898 453144
rect 254118 452548 254124 452600
rect 254176 452588 254182 452600
rect 282086 452588 282092 452600
rect 254176 452560 282092 452588
rect 254176 452548 254182 452560
rect 282086 452548 282092 452560
rect 282144 452548 282150 452600
rect 243170 452480 243176 452532
rect 243228 452520 243234 452532
rect 247034 452520 247040 452532
rect 243228 452492 247040 452520
rect 243228 452480 243234 452492
rect 247034 452480 247040 452492
rect 247092 452480 247098 452532
rect 255866 452480 255872 452532
rect 255924 452520 255930 452532
rect 284294 452520 284300 452532
rect 255924 452492 284300 452520
rect 255924 452480 255930 452492
rect 284294 452480 284300 452492
rect 284352 452480 284358 452532
rect 254578 452412 254584 452464
rect 254636 452452 254642 452464
rect 284386 452452 284392 452464
rect 254636 452424 284392 452452
rect 254636 452412 254642 452424
rect 284386 452412 284392 452424
rect 284444 452412 284450 452464
rect 253198 452344 253204 452396
rect 253256 452384 253262 452396
rect 284478 452384 284484 452396
rect 253256 452356 284484 452384
rect 253256 452344 253262 452356
rect 284478 452344 284484 452356
rect 284536 452344 284542 452396
rect 250714 452276 250720 452328
rect 250772 452316 250778 452328
rect 283006 452316 283012 452328
rect 250772 452288 283012 452316
rect 250772 452276 250778 452288
rect 283006 452276 283012 452288
rect 283064 452276 283070 452328
rect 251542 452208 251548 452260
rect 251600 452248 251606 452260
rect 284570 452248 284576 452260
rect 251600 452220 284576 452248
rect 251600 452208 251606 452220
rect 284570 452208 284576 452220
rect 284628 452208 284634 452260
rect 219710 452140 219716 452192
rect 219768 452180 219774 452192
rect 219986 452180 219992 452192
rect 219768 452152 219992 452180
rect 219768 452140 219774 452152
rect 219986 452140 219992 452152
rect 220044 452140 220050 452192
rect 248138 452140 248144 452192
rect 248196 452180 248202 452192
rect 281626 452180 281632 452192
rect 248196 452152 281632 452180
rect 248196 452140 248202 452152
rect 281626 452140 281632 452152
rect 281684 452140 281690 452192
rect 249426 452072 249432 452124
rect 249484 452112 249490 452124
rect 283098 452112 283104 452124
rect 249484 452084 283104 452112
rect 249484 452072 249490 452084
rect 283098 452072 283104 452084
rect 283156 452072 283162 452124
rect 245838 452004 245844 452056
rect 245896 452044 245902 452056
rect 280982 452044 280988 452056
rect 245896 452016 280988 452044
rect 245896 452004 245902 452016
rect 280982 452004 280988 452016
rect 281040 452004 281046 452056
rect 171778 451936 171784 451988
rect 171836 451976 171842 451988
rect 220722 451976 220728 451988
rect 171836 451948 220728 451976
rect 171836 451936 171842 451948
rect 220722 451936 220728 451948
rect 220780 451936 220786 451988
rect 234614 451936 234620 451988
rect 234672 451976 234678 451988
rect 235626 451976 235632 451988
rect 234672 451948 235632 451976
rect 234672 451936 234678 451948
rect 235626 451936 235632 451948
rect 235684 451936 235690 451988
rect 239030 451936 239036 451988
rect 239088 451976 239094 451988
rect 240042 451976 240048 451988
rect 239088 451948 240048 451976
rect 239088 451936 239094 451948
rect 240042 451936 240048 451948
rect 240100 451936 240106 451988
rect 241606 451936 241612 451988
rect 241664 451976 241670 451988
rect 242618 451976 242624 451988
rect 241664 451948 242624 451976
rect 241664 451936 241670 451948
rect 242618 451936 242624 451948
rect 242676 451936 242682 451988
rect 243078 451936 243084 451988
rect 243136 451976 243142 451988
rect 243906 451976 243912 451988
rect 243136 451948 243912 451976
rect 243136 451936 243142 451948
rect 243906 451936 243912 451948
rect 243964 451936 243970 451988
rect 247402 451936 247408 451988
rect 247460 451976 247466 451988
rect 299382 451976 299388 451988
rect 247460 451948 299388 451976
rect 247460 451936 247466 451948
rect 299382 451936 299388 451948
rect 299440 451936 299446 451988
rect 217318 451868 217324 451920
rect 217376 451908 217382 451920
rect 286318 451908 286324 451920
rect 217376 451880 286324 451908
rect 217376 451868 217382 451880
rect 286318 451868 286324 451880
rect 286376 451868 286382 451920
rect 214834 451256 214840 451308
rect 214892 451296 214898 451308
rect 221458 451296 221464 451308
rect 214892 451268 221464 451296
rect 214892 451256 214898 451268
rect 221458 451256 221464 451268
rect 221516 451256 221522 451308
rect 233970 451256 233976 451308
rect 234028 451296 234034 451308
rect 297818 451296 297824 451308
rect 234028 451268 297824 451296
rect 234028 451256 234034 451268
rect 297818 451256 297824 451268
rect 297876 451256 297882 451308
rect 229830 451188 229836 451240
rect 229888 451228 229894 451240
rect 242986 451228 242992 451240
rect 229888 451200 242992 451228
rect 229888 451188 229894 451200
rect 242986 451188 242992 451200
rect 243044 451228 243050 451240
rect 243538 451228 243544 451240
rect 243044 451200 243544 451228
rect 243044 451188 243050 451200
rect 243538 451188 243544 451200
rect 243596 451188 243602 451240
rect 189074 450916 189080 450968
rect 189132 450956 189138 450968
rect 230842 450956 230848 450968
rect 189132 450928 230848 450956
rect 189132 450916 189138 450928
rect 230842 450916 230848 450928
rect 230900 450916 230906 450968
rect 188430 450848 188436 450900
rect 188488 450888 188494 450900
rect 234246 450888 234252 450900
rect 188488 450860 234252 450888
rect 188488 450848 188494 450860
rect 234246 450848 234252 450860
rect 234304 450848 234310 450900
rect 187326 450780 187332 450832
rect 187384 450820 187390 450832
rect 233786 450820 233792 450832
rect 187384 450792 233792 450820
rect 187384 450780 187390 450792
rect 233786 450780 233792 450792
rect 233844 450780 233850 450832
rect 256050 450780 256056 450832
rect 256108 450820 256114 450832
rect 293218 450820 293224 450832
rect 256108 450792 293224 450820
rect 256108 450780 256114 450792
rect 293218 450780 293224 450792
rect 293276 450780 293282 450832
rect 187142 450712 187148 450764
rect 187200 450752 187206 450764
rect 233418 450752 233424 450764
rect 187200 450724 233424 450752
rect 187200 450712 187206 450724
rect 233418 450712 233424 450724
rect 233476 450712 233482 450764
rect 254762 450712 254768 450764
rect 254820 450752 254826 450764
rect 298002 450752 298008 450764
rect 254820 450724 298008 450752
rect 254820 450712 254826 450724
rect 298002 450712 298008 450724
rect 298060 450712 298066 450764
rect 187510 450644 187516 450696
rect 187568 450684 187574 450696
rect 234062 450684 234068 450696
rect 187568 450656 234068 450684
rect 187568 450644 187574 450656
rect 234062 450644 234068 450656
rect 234120 450644 234126 450696
rect 255682 450644 255688 450696
rect 255740 450684 255746 450696
rect 299750 450684 299756 450696
rect 255740 450656 299756 450684
rect 255740 450644 255746 450656
rect 299750 450644 299756 450656
rect 299808 450644 299814 450696
rect 187418 450576 187424 450628
rect 187476 450616 187482 450628
rect 255314 450616 255320 450628
rect 187476 450588 255320 450616
rect 187476 450576 187482 450588
rect 255314 450576 255320 450588
rect 255372 450576 255378 450628
rect 187234 450508 187240 450560
rect 187292 450548 187298 450560
rect 255406 450548 255412 450560
rect 187292 450520 255412 450548
rect 187292 450508 187298 450520
rect 255406 450508 255412 450520
rect 255464 450508 255470 450560
rect 3510 449828 3516 449880
rect 3568 449868 3574 449880
rect 223022 449868 223028 449880
rect 3568 449840 223028 449868
rect 3568 449828 3574 449840
rect 223022 449828 223028 449840
rect 223080 449828 223086 449880
rect 229738 449828 229744 449880
rect 229796 449868 229802 449880
rect 244918 449868 244924 449880
rect 229796 449840 244924 449868
rect 229796 449828 229802 449840
rect 244918 449828 244924 449840
rect 244976 449828 244982 449880
rect 204898 449760 204904 449812
rect 204956 449800 204962 449812
rect 232590 449800 232596 449812
rect 204956 449772 232596 449800
rect 204956 449760 204962 449772
rect 232590 449760 232596 449772
rect 232648 449760 232654 449812
rect 187050 449692 187056 449744
rect 187108 449732 187114 449744
rect 232774 449732 232780 449744
rect 187108 449704 232780 449732
rect 187108 449692 187114 449704
rect 232774 449692 232780 449704
rect 232832 449732 232838 449744
rect 238110 449732 238116 449744
rect 232832 449704 238116 449732
rect 232832 449692 232838 449704
rect 238110 449692 238116 449704
rect 238168 449692 238174 449744
rect 187602 449624 187608 449676
rect 187660 449664 187666 449676
rect 233050 449664 233056 449676
rect 187660 449636 233056 449664
rect 187660 449624 187666 449636
rect 233050 449624 233056 449636
rect 233108 449664 233114 449676
rect 239582 449664 239588 449676
rect 233108 449636 239588 449664
rect 233108 449624 233114 449636
rect 239582 449624 239588 449636
rect 239640 449624 239646 449676
rect 189994 449556 190000 449608
rect 190052 449596 190058 449608
rect 246114 449596 246120 449608
rect 190052 449568 246120 449596
rect 190052 449556 190058 449568
rect 246114 449556 246120 449568
rect 246172 449556 246178 449608
rect 253842 449556 253848 449608
rect 253900 449596 253906 449608
rect 281074 449596 281080 449608
rect 253900 449568 281080 449596
rect 253900 449556 253906 449568
rect 281074 449556 281080 449568
rect 281132 449556 281138 449608
rect 189902 449488 189908 449540
rect 189960 449528 189966 449540
rect 247310 449528 247316 449540
rect 189960 449500 247316 449528
rect 189960 449488 189966 449500
rect 247310 449488 247316 449500
rect 247368 449488 247374 449540
rect 252554 449488 252560 449540
rect 252612 449528 252618 449540
rect 281810 449528 281816 449540
rect 252612 449500 281816 449528
rect 252612 449488 252618 449500
rect 281810 449488 281816 449500
rect 281868 449488 281874 449540
rect 171870 449420 171876 449472
rect 171928 449460 171934 449472
rect 252370 449460 252376 449472
rect 171928 449432 252376 449460
rect 171928 449420 171934 449432
rect 252370 449420 252376 449432
rect 252428 449420 252434 449472
rect 281902 449460 281908 449472
rect 252480 449432 281908 449460
rect 140682 449352 140688 449404
rect 140740 449392 140746 449404
rect 244642 449392 244648 449404
rect 140740 449364 244648 449392
rect 140740 449352 140746 449364
rect 244642 449352 244648 449364
rect 244700 449352 244706 449404
rect 251266 449352 251272 449404
rect 251324 449392 251330 449404
rect 252480 449392 252508 449432
rect 281902 449420 281908 449432
rect 281960 449420 281966 449472
rect 281994 449392 282000 449404
rect 251324 449364 252508 449392
rect 252572 449364 282000 449392
rect 251324 449352 251330 449364
rect 115842 449284 115848 449336
rect 115900 449324 115906 449336
rect 238202 449324 238208 449336
rect 115900 449296 238208 449324
rect 115900 449284 115906 449296
rect 238202 449284 238208 449296
rect 238260 449284 238266 449336
rect 249886 449284 249892 449336
rect 249944 449324 249950 449336
rect 252572 449324 252600 449364
rect 281994 449352 282000 449364
rect 282052 449352 282058 449404
rect 249944 449296 252600 449324
rect 249944 449284 249950 449296
rect 252738 449284 252744 449336
rect 252796 449324 252802 449336
rect 281718 449324 281724 449336
rect 252796 449296 281724 449324
rect 252796 449284 252802 449296
rect 281718 449284 281724 449296
rect 281776 449284 281782 449336
rect 111702 449216 111708 449268
rect 111760 449256 111766 449268
rect 236914 449256 236920 449268
rect 111760 449228 236920 449256
rect 111760 449216 111766 449228
rect 236914 449216 236920 449228
rect 236972 449216 236978 449268
rect 246666 449216 246672 449268
rect 246724 449256 246730 449268
rect 298738 449256 298744 449268
rect 246724 449228 298744 449256
rect 246724 449216 246730 449228
rect 298738 449216 298744 449228
rect 298796 449216 298802 449268
rect 3878 449148 3884 449200
rect 3936 449188 3942 449200
rect 223114 449188 223120 449200
rect 3936 449160 223120 449188
rect 3936 449148 3942 449160
rect 223114 449148 223120 449160
rect 223172 449148 223178 449200
rect 241514 449148 241520 449200
rect 241572 449188 241578 449200
rect 298922 449188 298928 449200
rect 241572 449160 298928 449188
rect 241572 449148 241578 449160
rect 298922 449148 298928 449160
rect 298980 449148 298986 449200
rect 248690 449080 248696 449132
rect 248748 449120 248754 449132
rect 252738 449120 252744 449132
rect 248748 449092 252744 449120
rect 248748 449080 248754 449092
rect 252738 449080 252744 449092
rect 252796 449080 252802 449132
rect 255406 448944 255412 448996
rect 255464 448984 255470 448996
rect 293586 448984 293592 448996
rect 255464 448956 293592 448984
rect 255464 448944 255470 448956
rect 293586 448944 293592 448956
rect 293644 448944 293650 448996
rect 252186 448876 252192 448928
rect 252244 448916 252250 448928
rect 293678 448916 293684 448928
rect 252244 448888 293684 448916
rect 252244 448876 252250 448888
rect 293678 448876 293684 448888
rect 293736 448876 293742 448928
rect 249610 448808 249616 448860
rect 249668 448848 249674 448860
rect 293218 448848 293224 448860
rect 249668 448820 293224 448848
rect 249668 448808 249674 448820
rect 293218 448808 293224 448820
rect 293276 448808 293282 448860
rect 244274 448740 244280 448792
rect 244332 448780 244338 448792
rect 244918 448780 244924 448792
rect 244332 448752 244924 448780
rect 244332 448740 244338 448752
rect 244918 448740 244924 448752
rect 244976 448740 244982 448792
rect 247034 448740 247040 448792
rect 247092 448780 247098 448792
rect 293862 448780 293868 448792
rect 247092 448752 293868 448780
rect 247092 448740 247098 448752
rect 293862 448740 293868 448752
rect 293920 448740 293926 448792
rect 244090 448672 244096 448724
rect 244148 448712 244154 448724
rect 296530 448712 296536 448724
rect 244148 448684 296536 448712
rect 244148 448672 244154 448684
rect 296530 448672 296536 448684
rect 296588 448672 296594 448724
rect 230474 448604 230480 448656
rect 230532 448644 230538 448656
rect 293402 448644 293408 448656
rect 230532 448616 293408 448644
rect 230532 448604 230538 448616
rect 293402 448604 293408 448616
rect 293460 448604 293466 448656
rect 230290 448536 230296 448588
rect 230348 448576 230354 448588
rect 293770 448576 293776 448588
rect 230348 448548 293776 448576
rect 230348 448536 230354 448548
rect 293770 448536 293776 448548
rect 293828 448536 293834 448588
rect 23474 448468 23480 448520
rect 23532 448508 23538 448520
rect 222194 448508 222200 448520
rect 23532 448480 222200 448508
rect 23532 448468 23538 448480
rect 222194 448468 222200 448480
rect 222252 448508 222258 448520
rect 222930 448508 222936 448520
rect 222252 448480 222936 448508
rect 222252 448468 222258 448480
rect 222930 448468 222936 448480
rect 222988 448468 222994 448520
rect 238110 448468 238116 448520
rect 238168 448508 238174 448520
rect 297634 448508 297640 448520
rect 238168 448480 297640 448508
rect 238168 448468 238174 448480
rect 297634 448468 297640 448480
rect 297692 448468 297698 448520
rect 239582 448400 239588 448452
rect 239640 448440 239646 448452
rect 297726 448440 297732 448452
rect 239640 448412 297732 448440
rect 239640 448400 239646 448412
rect 297726 448400 297732 448412
rect 297784 448400 297790 448452
rect 222838 448332 222844 448384
rect 222896 448372 222902 448384
rect 231946 448372 231952 448384
rect 222896 448344 231952 448372
rect 222896 448332 222902 448344
rect 231946 448332 231952 448344
rect 232004 448372 232010 448384
rect 232498 448372 232504 448384
rect 232004 448344 232504 448372
rect 232004 448332 232010 448344
rect 232498 448332 232504 448344
rect 232556 448332 232562 448384
rect 297910 448372 297916 448384
rect 244246 448344 297916 448372
rect 233418 448264 233424 448316
rect 233476 448304 233482 448316
rect 244246 448304 244274 448344
rect 297910 448332 297916 448344
rect 297968 448332 297974 448384
rect 297450 448304 297456 448316
rect 233476 448276 244274 448304
rect 248386 448276 297456 448304
rect 233476 448264 233482 448276
rect 184198 448196 184204 448248
rect 184256 448236 184262 448248
rect 221642 448236 221648 448248
rect 184256 448208 221648 448236
rect 184256 448196 184262 448208
rect 221642 448196 221648 448208
rect 221700 448196 221706 448248
rect 226978 448196 226984 448248
rect 227036 448236 227042 448248
rect 240410 448236 240416 448248
rect 227036 448208 240416 448236
rect 227036 448196 227042 448208
rect 240410 448196 240416 448208
rect 240468 448196 240474 448248
rect 3970 448128 3976 448180
rect 4028 448168 4034 448180
rect 223482 448168 223488 448180
rect 4028 448140 223488 448168
rect 4028 448128 4034 448140
rect 223482 448128 223488 448140
rect 223540 448128 223546 448180
rect 233786 448128 233792 448180
rect 233844 448168 233850 448180
rect 248386 448168 248414 448276
rect 297450 448264 297456 448276
rect 297508 448264 297514 448316
rect 255314 448196 255320 448248
rect 255372 448236 255378 448248
rect 256234 448236 256240 448248
rect 255372 448208 256240 448236
rect 255372 448196 255378 448208
rect 256234 448196 256240 448208
rect 256292 448236 256298 448248
rect 297542 448236 297548 448248
rect 256292 448208 297548 448236
rect 256292 448196 256298 448208
rect 297542 448196 297548 448208
rect 297600 448196 297606 448248
rect 233844 448140 248414 448168
rect 233844 448128 233850 448140
rect 3694 448060 3700 448112
rect 3752 448100 3758 448112
rect 222930 448100 222936 448112
rect 3752 448072 222936 448100
rect 3752 448060 3758 448072
rect 222930 448060 222936 448072
rect 222988 448060 222994 448112
rect 3602 447992 3608 448044
rect 3660 448032 3666 448044
rect 222562 448032 222568 448044
rect 3660 448004 222568 448032
rect 3660 447992 3666 448004
rect 222562 447992 222568 448004
rect 222620 447992 222626 448044
rect 3786 447924 3792 447976
rect 3844 447964 3850 447976
rect 223298 447964 223304 447976
rect 3844 447936 223304 447964
rect 3844 447924 3850 447936
rect 223298 447924 223304 447936
rect 223356 447924 223362 447976
rect 231762 447924 231768 447976
rect 231820 447964 231826 447976
rect 239674 447964 239680 447976
rect 231820 447936 239680 447964
rect 231820 447924 231826 447936
rect 239674 447924 239680 447936
rect 239732 447924 239738 447976
rect 3418 447856 3424 447908
rect 3476 447896 3482 447908
rect 222378 447896 222384 447908
rect 3476 447868 222384 447896
rect 3476 447856 3482 447868
rect 222378 447856 222384 447868
rect 222436 447856 222442 447908
rect 236730 447856 236736 447908
rect 236788 447896 236794 447908
rect 253290 447896 253296 447908
rect 236788 447868 253296 447896
rect 236788 447856 236794 447868
rect 253290 447856 253296 447868
rect 253348 447856 253354 447908
rect 3234 447788 3240 447840
rect 3292 447828 3298 447840
rect 224770 447828 224776 447840
rect 3292 447800 224776 447828
rect 3292 447788 3298 447800
rect 224770 447788 224776 447800
rect 224828 447788 224834 447840
rect 226242 447788 226248 447840
rect 226300 447828 226306 447840
rect 238386 447828 238392 447840
rect 226300 447800 238392 447828
rect 226300 447788 226306 447800
rect 238386 447788 238392 447800
rect 238444 447788 238450 447840
rect 245746 447788 245752 447840
rect 245804 447828 245810 447840
rect 296070 447828 296076 447840
rect 245804 447800 296076 447828
rect 245804 447788 245810 447800
rect 296070 447788 296076 447800
rect 296128 447788 296134 447840
rect 246206 447720 246212 447772
rect 246264 447760 246270 447772
rect 246482 447760 246488 447772
rect 246264 447732 246488 447760
rect 246264 447720 246270 447732
rect 246482 447720 246488 447732
rect 246540 447720 246546 447772
rect 244734 447652 244740 447704
rect 244792 447692 244798 447704
rect 249978 447692 249984 447704
rect 244792 447664 249984 447692
rect 244792 447652 244798 447664
rect 249978 447652 249984 447664
rect 250036 447652 250042 447704
rect 240594 447584 240600 447636
rect 240652 447624 240658 447636
rect 240652 447596 248414 447624
rect 240652 447584 240658 447596
rect 230106 447516 230112 447568
rect 230164 447556 230170 447568
rect 230164 447528 235396 447556
rect 230164 447516 230170 447528
rect 219434 447380 219440 447432
rect 219492 447420 219498 447432
rect 219894 447420 219900 447432
rect 219492 447392 219900 447420
rect 219492 447380 219498 447392
rect 219894 447380 219900 447392
rect 219952 447380 219958 447432
rect 231762 447380 231768 447432
rect 231820 447420 231826 447432
rect 231820 447392 234614 447420
rect 231820 447380 231826 447392
rect 214006 447312 214012 447364
rect 214064 447352 214070 447364
rect 215018 447352 215024 447364
rect 214064 447324 215024 447352
rect 214064 447312 214070 447324
rect 215018 447312 215024 447324
rect 215076 447312 215082 447364
rect 215294 447312 215300 447364
rect 215352 447352 215358 447364
rect 216122 447352 216128 447364
rect 215352 447324 216128 447352
rect 215352 447312 215358 447324
rect 216122 447312 216128 447324
rect 216180 447312 216186 447364
rect 217134 447312 217140 447364
rect 217192 447352 217198 447364
rect 217594 447352 217600 447364
rect 217192 447324 217600 447352
rect 217192 447312 217198 447324
rect 217594 447312 217600 447324
rect 217652 447312 217658 447364
rect 218054 447312 218060 447364
rect 218112 447352 218118 447364
rect 218882 447352 218888 447364
rect 218112 447324 218888 447352
rect 218112 447312 218118 447324
rect 218882 447312 218888 447324
rect 218940 447312 218946 447364
rect 220998 447312 221004 447364
rect 221056 447352 221062 447364
rect 221826 447352 221832 447364
rect 221056 447324 221832 447352
rect 221056 447312 221062 447324
rect 221826 447312 221832 447324
rect 221884 447312 221890 447364
rect 214190 447244 214196 447296
rect 214248 447284 214254 447296
rect 215202 447284 215208 447296
rect 214248 447256 215208 447284
rect 214248 447244 214254 447256
rect 215202 447244 215208 447256
rect 215260 447244 215266 447296
rect 215846 447244 215852 447296
rect 215904 447284 215910 447296
rect 216306 447284 216312 447296
rect 215904 447256 216312 447284
rect 215904 447244 215910 447256
rect 216306 447244 216312 447256
rect 216364 447244 216370 447296
rect 216766 447244 216772 447296
rect 216824 447284 216830 447296
rect 217778 447284 217784 447296
rect 216824 447256 217784 447284
rect 216824 447244 216830 447256
rect 217778 447244 217784 447256
rect 217836 447244 217842 447296
rect 218606 447244 218612 447296
rect 218664 447284 218670 447296
rect 219250 447284 219256 447296
rect 218664 447256 219256 447284
rect 218664 447244 218670 447256
rect 219250 447244 219256 447256
rect 219308 447244 219314 447296
rect 220906 447244 220912 447296
rect 220964 447284 220970 447296
rect 221366 447284 221372 447296
rect 220964 447256 221372 447284
rect 220964 447244 220970 447256
rect 221366 447244 221372 447256
rect 221424 447244 221430 447296
rect 224218 447244 224224 447296
rect 224276 447284 224282 447296
rect 224678 447284 224684 447296
rect 224276 447256 224684 447284
rect 224276 447244 224282 447256
rect 224678 447244 224684 447256
rect 224736 447244 224742 447296
rect 234586 447284 234614 447392
rect 235368 447352 235396 447528
rect 241882 447516 241888 447568
rect 241940 447556 241946 447568
rect 246298 447556 246304 447568
rect 241940 447528 246304 447556
rect 241940 447516 241946 447528
rect 246298 447516 246304 447528
rect 246356 447516 246362 447568
rect 244366 447448 244372 447500
rect 244424 447488 244430 447500
rect 245562 447488 245568 447500
rect 244424 447460 245568 447488
rect 244424 447448 244430 447460
rect 245562 447448 245568 447460
rect 245620 447448 245626 447500
rect 245838 447448 245844 447500
rect 245896 447488 245902 447500
rect 246850 447488 246856 447500
rect 245896 447460 246856 447488
rect 245896 447448 245902 447460
rect 246850 447448 246856 447460
rect 246908 447448 246914 447500
rect 248386 447488 248414 447596
rect 251358 447516 251364 447568
rect 251416 447556 251422 447568
rect 251818 447556 251824 447568
rect 251416 447528 251824 447556
rect 251416 447516 251422 447528
rect 251818 447516 251824 447528
rect 251876 447516 251882 447568
rect 298002 447488 298008 447500
rect 248386 447460 298008 447488
rect 298002 447448 298008 447460
rect 298060 447448 298066 447500
rect 235442 447380 235448 447432
rect 235500 447420 235506 447432
rect 293494 447420 293500 447432
rect 235500 447392 293500 447420
rect 235500 447380 235506 447392
rect 293494 447380 293500 447392
rect 293552 447380 293558 447432
rect 293126 447352 293132 447364
rect 235368 447324 293132 447352
rect 293126 447312 293132 447324
rect 293184 447312 293190 447364
rect 296622 447284 296628 447296
rect 234586 447256 296628 447284
rect 296622 447244 296628 447256
rect 296680 447244 296686 447296
rect 220814 447176 220820 447228
rect 220872 447216 220878 447228
rect 222010 447216 222016 447228
rect 220872 447188 222016 447216
rect 220872 447176 220878 447188
rect 222010 447176 222016 447188
rect 222068 447176 222074 447228
rect 223298 447176 223304 447228
rect 223356 447216 223362 447228
rect 298646 447216 298652 447228
rect 223356 447188 298652 447216
rect 223356 447176 223362 447188
rect 298646 447176 298652 447188
rect 298704 447176 298710 447228
rect 213362 447108 213368 447160
rect 213420 447148 213426 447160
rect 296254 447148 296260 447160
rect 213420 447120 296260 447148
rect 213420 447108 213426 447120
rect 296254 447108 296260 447120
rect 296312 447108 296318 447160
rect 229922 447040 229928 447092
rect 229980 447080 229986 447092
rect 230658 447080 230664 447092
rect 229980 447052 230664 447080
rect 229980 447040 229986 447052
rect 230658 447040 230664 447052
rect 230716 447040 230722 447092
rect 243722 447040 243728 447092
rect 243780 447080 243786 447092
rect 246206 447080 246212 447092
rect 243780 447052 246212 447080
rect 243780 447040 243786 447052
rect 246206 447040 246212 447052
rect 246264 447040 246270 447092
rect 282270 447080 282276 447092
rect 253906 447052 282276 447080
rect 250346 446972 250352 447024
rect 250404 447012 250410 447024
rect 253906 447012 253934 447052
rect 282270 447040 282276 447052
rect 282328 447040 282334 447092
rect 283558 447012 283564 447024
rect 250404 446984 253934 447012
rect 258736 446984 283564 447012
rect 250404 446972 250410 446984
rect 247770 446904 247776 446956
rect 247828 446944 247834 446956
rect 258534 446944 258540 446956
rect 247828 446916 258540 446944
rect 247828 446904 247834 446916
rect 258534 446904 258540 446916
rect 258592 446904 258598 446956
rect 250162 446836 250168 446888
rect 250220 446876 250226 446888
rect 258736 446876 258764 446984
rect 283558 446972 283564 446984
rect 283616 446972 283622 447024
rect 258902 446904 258908 446956
rect 258960 446944 258966 446956
rect 282178 446944 282184 446956
rect 258960 446916 282184 446944
rect 258960 446904 258966 446916
rect 282178 446904 282184 446916
rect 282236 446904 282242 446956
rect 250220 446848 258764 446876
rect 250220 446836 250226 446848
rect 258810 446836 258816 446888
rect 258868 446876 258874 446888
rect 285030 446876 285036 446888
rect 258868 446848 285036 446876
rect 258868 446836 258874 446848
rect 285030 446836 285036 446848
rect 285088 446836 285094 446888
rect 224954 446768 224960 446820
rect 225012 446808 225018 446820
rect 225598 446808 225604 446820
rect 225012 446780 225604 446808
rect 225012 446768 225018 446780
rect 225598 446768 225604 446780
rect 225656 446808 225662 446820
rect 248966 446808 248972 446820
rect 225656 446780 248972 446808
rect 225656 446768 225662 446780
rect 248966 446768 248972 446780
rect 249024 446768 249030 446820
rect 251450 446768 251456 446820
rect 251508 446808 251514 446820
rect 289170 446808 289176 446820
rect 251508 446780 289176 446808
rect 251508 446768 251514 446780
rect 289170 446768 289176 446780
rect 289228 446768 289234 446820
rect 4982 446700 4988 446752
rect 5040 446740 5046 446752
rect 227714 446740 227720 446752
rect 5040 446712 227720 446740
rect 5040 446700 5046 446712
rect 227714 446700 227720 446712
rect 227772 446700 227778 446752
rect 252738 446700 252744 446752
rect 252796 446740 252802 446752
rect 293310 446740 293316 446752
rect 252796 446712 293316 446740
rect 252796 446700 252802 446712
rect 293310 446700 293316 446712
rect 293368 446700 293374 446752
rect 4798 446632 4804 446684
rect 4856 446672 4862 446684
rect 228818 446672 228824 446684
rect 4856 446644 228824 446672
rect 4856 446632 4862 446644
rect 228818 446632 228824 446644
rect 228876 446632 228882 446684
rect 246390 446632 246396 446684
rect 246448 446672 246454 446684
rect 287698 446672 287704 446684
rect 246448 446644 287704 446672
rect 246448 446632 246454 446644
rect 287698 446632 287704 446644
rect 287756 446632 287762 446684
rect 3510 446564 3516 446616
rect 3568 446604 3574 446616
rect 229370 446604 229376 446616
rect 3568 446576 229376 446604
rect 3568 446564 3574 446576
rect 229370 446564 229376 446576
rect 229428 446564 229434 446616
rect 247586 446564 247592 446616
rect 247644 446604 247650 446616
rect 289078 446604 289084 446616
rect 247644 446576 289084 446604
rect 247644 446564 247650 446576
rect 289078 446564 289084 446576
rect 289136 446564 289142 446616
rect 188982 446496 188988 446548
rect 189040 446536 189046 446548
rect 220538 446536 220544 446548
rect 189040 446508 220544 446536
rect 189040 446496 189046 446508
rect 220538 446496 220544 446508
rect 220596 446496 220602 446548
rect 238110 446496 238116 446548
rect 238168 446536 238174 446548
rect 255406 446536 255412 446548
rect 238168 446508 255412 446536
rect 238168 446496 238174 446508
rect 255406 446496 255412 446508
rect 255464 446496 255470 446548
rect 256602 446496 256608 446548
rect 256660 446536 256666 446548
rect 298094 446536 298100 446548
rect 256660 446508 298100 446536
rect 256660 446496 256666 446508
rect 298094 446496 298100 446508
rect 298152 446496 298158 446548
rect 188890 446428 188896 446480
rect 188948 446468 188954 446480
rect 220354 446468 220360 446480
rect 188948 446440 220360 446468
rect 188948 446428 188954 446440
rect 220354 446428 220360 446440
rect 220412 446428 220418 446480
rect 233234 446428 233240 446480
rect 233292 446468 233298 446480
rect 251726 446468 251732 446480
rect 233292 446440 251732 446468
rect 233292 446428 233298 446440
rect 251726 446428 251732 446440
rect 251784 446428 251790 446480
rect 256510 446428 256516 446480
rect 256568 446468 256574 446480
rect 299842 446468 299848 446480
rect 256568 446440 299848 446468
rect 256568 446428 256574 446440
rect 299842 446428 299848 446440
rect 299900 446428 299906 446480
rect 172054 446360 172060 446412
rect 172112 446400 172118 446412
rect 245930 446400 245936 446412
rect 172112 446372 245936 446400
rect 172112 446360 172118 446372
rect 245930 446360 245936 446372
rect 245988 446360 245994 446412
rect 253934 446360 253940 446412
rect 253992 446400 253998 446412
rect 298830 446400 298836 446412
rect 253992 446372 298836 446400
rect 253992 446360 253998 446372
rect 298830 446360 298836 446372
rect 298888 446360 298894 446412
rect 3602 446292 3608 446344
rect 3660 446332 3666 446344
rect 228634 446332 228640 446344
rect 3660 446304 228640 446332
rect 3660 446292 3666 446304
rect 228634 446292 228640 446304
rect 228692 446292 228698 446344
rect 255314 446292 255320 446344
rect 255372 446332 255378 446344
rect 286410 446332 286416 446344
rect 255372 446304 286416 446332
rect 255372 446292 255378 446304
rect 286410 446292 286416 446304
rect 286468 446292 286474 446344
rect 209130 446224 209136 446276
rect 209188 446264 209194 446276
rect 230382 446264 230388 446276
rect 209188 446236 230388 446264
rect 209188 446224 209194 446236
rect 230382 446224 230388 446236
rect 230440 446224 230446 446276
rect 252922 446224 252928 446276
rect 252980 446264 252986 446276
rect 282362 446264 282368 446276
rect 252980 446236 282368 446264
rect 252980 446224 252986 446236
rect 282362 446224 282368 446236
rect 282420 446224 282426 446276
rect 221642 446156 221648 446208
rect 221700 446196 221706 446208
rect 246942 446196 246948 446208
rect 221700 446168 246948 446196
rect 221700 446156 221706 446168
rect 246942 446156 246948 446168
rect 247000 446156 247006 446208
rect 248874 446156 248880 446208
rect 248932 446196 248938 446208
rect 258810 446196 258816 446208
rect 248932 446168 258816 446196
rect 248932 446156 248938 446168
rect 258810 446156 258816 446168
rect 258868 446156 258874 446208
rect 5166 446088 5172 446140
rect 5224 446128 5230 446140
rect 226058 446128 226064 446140
rect 5224 446100 226064 446128
rect 5224 446088 5230 446100
rect 226058 446088 226064 446100
rect 226116 446088 226122 446140
rect 234338 446088 234344 446140
rect 234396 446128 234402 446140
rect 256326 446128 256332 446140
rect 234396 446100 256332 446128
rect 234396 446088 234402 446100
rect 256326 446088 256332 446100
rect 256384 446088 256390 446140
rect 5074 446020 5080 446072
rect 5132 446060 5138 446072
rect 226610 446060 226616 446072
rect 5132 446032 226616 446060
rect 5132 446020 5138 446032
rect 226610 446020 226616 446032
rect 226668 446020 226674 446072
rect 216582 445952 216588 446004
rect 216640 445992 216646 446004
rect 225506 445992 225512 446004
rect 216640 445964 225512 445992
rect 216640 445952 216646 445964
rect 225506 445952 225512 445964
rect 225564 445952 225570 446004
rect 249886 445992 249892 446004
rect 241486 445964 249892 445992
rect 213822 445884 213828 445936
rect 213880 445924 213886 445936
rect 228082 445924 228088 445936
rect 213880 445896 228088 445924
rect 213880 445884 213886 445896
rect 228082 445884 228088 445896
rect 228140 445884 228146 445936
rect 211062 445816 211068 445868
rect 211120 445856 211126 445868
rect 226978 445856 226984 445868
rect 211120 445828 226984 445856
rect 211120 445816 211126 445828
rect 226978 445816 226984 445828
rect 227036 445816 227042 445868
rect 232866 445816 232872 445868
rect 232924 445856 232930 445868
rect 241486 445856 241514 445964
rect 249886 445952 249892 445964
rect 249944 445952 249950 446004
rect 245378 445884 245384 445936
rect 245436 445924 245442 445936
rect 245436 445896 246528 445924
rect 245436 445884 245442 445896
rect 232924 445828 241514 445856
rect 232924 445816 232930 445828
rect 245010 445816 245016 445868
rect 245068 445856 245074 445868
rect 246298 445856 246304 445868
rect 245068 445828 246304 445856
rect 245068 445816 245074 445828
rect 246298 445816 246304 445828
rect 246356 445816 246362 445868
rect 246500 445856 246528 445896
rect 256510 445856 256516 445868
rect 246500 445828 256516 445856
rect 256510 445816 256516 445828
rect 256568 445816 256574 445868
rect 208394 445748 208400 445800
rect 208452 445788 208458 445800
rect 227530 445788 227536 445800
rect 208452 445760 227536 445788
rect 208452 445748 208458 445760
rect 227530 445748 227536 445760
rect 227588 445748 227594 445800
rect 235994 445748 236000 445800
rect 236052 445788 236058 445800
rect 238018 445788 238024 445800
rect 236052 445760 238024 445788
rect 236052 445748 236058 445760
rect 238018 445748 238024 445760
rect 238076 445748 238082 445800
rect 240226 445748 240232 445800
rect 240284 445788 240290 445800
rect 295886 445788 295892 445800
rect 240284 445760 295892 445788
rect 240284 445748 240290 445760
rect 295886 445748 295892 445760
rect 295944 445748 295950 445800
rect 227898 445680 227904 445732
rect 227956 445720 227962 445732
rect 228450 445720 228456 445732
rect 227956 445692 228456 445720
rect 227956 445680 227962 445692
rect 228450 445680 228456 445692
rect 228508 445680 228514 445732
rect 196618 445544 196624 445596
rect 196676 445584 196682 445596
rect 227898 445584 227904 445596
rect 196676 445556 227904 445584
rect 196676 445544 196682 445556
rect 227898 445544 227904 445556
rect 227956 445544 227962 445596
rect 225506 445476 225512 445528
rect 225564 445516 225570 445528
rect 266170 445516 266176 445528
rect 225564 445488 266176 445516
rect 225564 445476 225570 445488
rect 266170 445476 266176 445488
rect 266228 445476 266234 445528
rect 199654 445408 199660 445460
rect 199712 445448 199718 445460
rect 226242 445448 226248 445460
rect 199712 445420 226248 445448
rect 199712 445408 199718 445420
rect 226242 445408 226248 445420
rect 226300 445408 226306 445460
rect 196710 445340 196716 445392
rect 196768 445380 196774 445392
rect 226794 445380 226800 445392
rect 196768 445352 226800 445380
rect 196768 445340 196774 445352
rect 226794 445340 226800 445352
rect 226852 445340 226858 445392
rect 254118 445340 254124 445392
rect 254176 445380 254182 445392
rect 255130 445380 255136 445392
rect 254176 445352 255136 445380
rect 254176 445340 254182 445352
rect 255130 445340 255136 445352
rect 255188 445340 255194 445392
rect 210786 445272 210792 445324
rect 210844 445312 210850 445324
rect 273898 445312 273904 445324
rect 210844 445284 273904 445312
rect 210844 445272 210850 445284
rect 273898 445272 273904 445284
rect 273956 445272 273962 445324
rect 199562 445204 199568 445256
rect 199620 445244 199626 445256
rect 227346 445244 227352 445256
rect 199620 445216 227352 445244
rect 199620 445204 199626 445216
rect 227346 445204 227352 445216
rect 227404 445204 227410 445256
rect 236270 445204 236276 445256
rect 236328 445244 236334 445256
rect 237282 445244 237288 445256
rect 236328 445216 237288 445244
rect 236328 445204 236334 445216
rect 237282 445204 237288 445216
rect 237340 445204 237346 445256
rect 237926 445204 237932 445256
rect 237984 445244 237990 445256
rect 238570 445244 238576 445256
rect 237984 445216 238576 445244
rect 237984 445204 237990 445216
rect 238570 445204 238576 445216
rect 238628 445204 238634 445256
rect 238846 445204 238852 445256
rect 238904 445244 238910 445256
rect 239858 445244 239864 445256
rect 238904 445216 239864 445244
rect 238904 445204 238910 445216
rect 239858 445204 239864 445216
rect 239916 445204 239922 445256
rect 240318 445204 240324 445256
rect 240376 445244 240382 445256
rect 241330 445244 241336 445256
rect 240376 445216 241336 445244
rect 240376 445204 240382 445216
rect 241330 445204 241336 445216
rect 241388 445204 241394 445256
rect 241790 445204 241796 445256
rect 241848 445244 241854 445256
rect 242434 445244 242440 445256
rect 241848 445216 242440 445244
rect 241848 445204 241854 445216
rect 242434 445204 242440 445216
rect 242492 445204 242498 445256
rect 247126 445204 247132 445256
rect 247184 445244 247190 445256
rect 248322 445244 248328 445256
rect 247184 445216 248328 445244
rect 247184 445204 247190 445216
rect 248322 445204 248328 445216
rect 248380 445204 248386 445256
rect 248414 445204 248420 445256
rect 248472 445244 248478 445256
rect 249058 445244 249064 445256
rect 248472 445216 249064 445244
rect 248472 445204 248478 445216
rect 249058 445204 249064 445216
rect 249116 445204 249122 445256
rect 3786 445136 3792 445188
rect 3844 445176 3850 445188
rect 208394 445176 208400 445188
rect 3844 445148 208400 445176
rect 3844 445136 3850 445148
rect 208394 445136 208400 445148
rect 208452 445136 208458 445188
rect 213546 445136 213552 445188
rect 213604 445176 213610 445188
rect 269850 445176 269856 445188
rect 213604 445148 269856 445176
rect 213604 445136 213610 445148
rect 269850 445136 269856 445148
rect 269908 445136 269914 445188
rect 3878 445068 3884 445120
rect 3936 445108 3942 445120
rect 211062 445108 211068 445120
rect 3936 445080 211068 445108
rect 3936 445068 3942 445080
rect 211062 445068 211068 445080
rect 211120 445068 211126 445120
rect 215662 445068 215668 445120
rect 215720 445108 215726 445120
rect 216490 445108 216496 445120
rect 215720 445080 216496 445108
rect 215720 445068 215726 445080
rect 216490 445068 216496 445080
rect 216548 445068 216554 445120
rect 217042 445068 217048 445120
rect 217100 445108 217106 445120
rect 217318 445108 217324 445120
rect 217100 445080 217324 445108
rect 217100 445068 217106 445080
rect 217318 445068 217324 445080
rect 217376 445068 217382 445120
rect 218238 445068 218244 445120
rect 218296 445108 218302 445120
rect 218698 445108 218704 445120
rect 218296 445080 218704 445108
rect 218296 445068 218302 445080
rect 218698 445068 218704 445080
rect 218756 445068 218762 445120
rect 229554 445068 229560 445120
rect 229612 445108 229618 445120
rect 268470 445108 268476 445120
rect 229612 445080 268476 445108
rect 229612 445068 229618 445080
rect 268470 445068 268476 445080
rect 268528 445068 268534 445120
rect 3694 445000 3700 445052
rect 3752 445040 3758 445052
rect 213822 445040 213828 445052
rect 3752 445012 213828 445040
rect 3752 445000 3758 445012
rect 213822 445000 213828 445012
rect 213880 445000 213886 445052
rect 246942 445000 246948 445052
rect 247000 445040 247006 445052
rect 299474 445040 299480 445052
rect 247000 445012 299480 445040
rect 247000 445000 247006 445012
rect 299474 445000 299480 445012
rect 299532 445000 299538 445052
rect 226794 444932 226800 444984
rect 226852 444972 226858 444984
rect 267090 444972 267096 444984
rect 226852 444944 267096 444972
rect 226852 444932 226858 444944
rect 267090 444932 267096 444944
rect 267148 444932 267154 444984
rect 199470 444864 199476 444916
rect 199528 444904 199534 444916
rect 228450 444904 228456 444916
rect 199528 444876 228456 444904
rect 199528 444864 199534 444876
rect 228450 444864 228456 444876
rect 228508 444864 228514 444916
rect 212442 444796 212448 444848
rect 212500 444836 212506 444848
rect 268378 444836 268384 444848
rect 212500 444808 268384 444836
rect 212500 444796 212506 444808
rect 268378 444796 268384 444808
rect 268436 444796 268442 444848
rect 211338 444728 211344 444780
rect 211396 444768 211402 444780
rect 275278 444768 275284 444780
rect 211396 444740 275284 444768
rect 211396 444728 211402 444740
rect 275278 444728 275284 444740
rect 275336 444728 275342 444780
rect 210970 444660 210976 444712
rect 211028 444700 211034 444712
rect 278038 444700 278044 444712
rect 211028 444672 278044 444700
rect 211028 444660 211034 444672
rect 278038 444660 278044 444672
rect 278096 444660 278102 444712
rect 213914 444592 213920 444644
rect 213972 444632 213978 444644
rect 296438 444632 296444 444644
rect 213972 444604 296444 444632
rect 213972 444592 213978 444604
rect 296438 444592 296444 444604
rect 296496 444592 296502 444644
rect 213730 444524 213736 444576
rect 213788 444564 213794 444576
rect 299290 444564 299296 444576
rect 213788 444536 299296 444564
rect 213788 444524 213794 444536
rect 299290 444524 299296 444536
rect 299348 444524 299354 444576
rect 98638 444456 98644 444508
rect 98696 444496 98702 444508
rect 225690 444496 225696 444508
rect 98696 444468 225696 444496
rect 98696 444456 98702 444468
rect 225690 444456 225696 444468
rect 225748 444456 225754 444508
rect 253474 444456 253480 444508
rect 253532 444496 253538 444508
rect 293310 444496 293316 444508
rect 253532 444468 293316 444496
rect 253532 444456 253538 444468
rect 293310 444456 293316 444468
rect 293368 444456 293374 444508
rect 13078 444388 13084 444440
rect 13136 444428 13142 444440
rect 225138 444428 225144 444440
rect 13136 444400 225144 444428
rect 13136 444388 13142 444400
rect 225138 444388 225144 444400
rect 225196 444388 225202 444440
rect 254394 444388 254400 444440
rect 254452 444428 254458 444440
rect 266078 444428 266084 444440
rect 254452 444400 266084 444428
rect 254452 444388 254458 444400
rect 266078 444388 266084 444400
rect 266136 444388 266142 444440
rect 251542 444184 251548 444236
rect 251600 444224 251606 444236
rect 252002 444224 252008 444236
rect 251600 444196 252008 444224
rect 251600 444184 251606 444196
rect 252002 444184 252008 444196
rect 252060 444184 252066 444236
rect 212994 444048 213000 444100
rect 213052 444088 213058 444100
rect 220262 444088 220268 444100
rect 213052 444060 220268 444088
rect 213052 444048 213058 444060
rect 220262 444048 220268 444060
rect 220320 444048 220326 444100
rect 256510 443844 256516 443896
rect 256568 443884 256574 443896
rect 295794 443884 295800 443896
rect 256568 443856 295800 443884
rect 256568 443844 256574 443856
rect 295794 443844 295800 443856
rect 295852 443844 295858 443896
rect 214190 443776 214196 443828
rect 214248 443816 214254 443828
rect 217502 443816 217508 443828
rect 214248 443788 217508 443816
rect 214248 443776 214254 443788
rect 217502 443776 217508 443788
rect 217560 443776 217566 443828
rect 254486 443776 254492 443828
rect 254544 443816 254550 443828
rect 256142 443816 256148 443828
rect 254544 443788 256148 443816
rect 254544 443776 254550 443788
rect 256142 443776 256148 443788
rect 256200 443776 256206 443828
rect 256326 443776 256332 443828
rect 256384 443816 256390 443828
rect 297358 443816 297364 443828
rect 256384 443788 297364 443816
rect 256384 443776 256390 443788
rect 297358 443776 297364 443788
rect 297416 443776 297422 443828
rect 249886 443708 249892 443760
rect 249944 443748 249950 443760
rect 297450 443748 297456 443760
rect 249944 443720 297456 443748
rect 249944 443708 249950 443720
rect 297450 443708 297456 443720
rect 297508 443708 297514 443760
rect 3234 443640 3240 443692
rect 3292 443680 3298 443692
rect 216582 443680 216588 443692
rect 3292 443652 216588 443680
rect 3292 443640 3298 443652
rect 216582 443640 216588 443652
rect 216640 443640 216646 443692
rect 229830 443680 229836 443692
rect 222166 443652 229836 443680
rect 212534 443572 212540 443624
rect 212592 443612 212598 443624
rect 222166 443612 222194 443652
rect 229830 443640 229836 443652
rect 229888 443640 229894 443692
rect 234430 443640 234436 443692
rect 234488 443680 234494 443692
rect 239950 443680 239956 443692
rect 234488 443652 239956 443680
rect 234488 443640 234494 443652
rect 239950 443640 239956 443652
rect 240008 443640 240014 443692
rect 242710 443680 242716 443692
rect 240106 443652 242716 443680
rect 212592 443584 222194 443612
rect 224926 443584 234614 443612
rect 212592 443572 212598 443584
rect 213748 443516 216444 443544
rect 199378 443436 199384 443488
rect 199436 443476 199442 443488
rect 212534 443476 212540 443488
rect 199436 443448 212540 443476
rect 199436 443436 199442 443448
rect 212534 443436 212540 443448
rect 212592 443436 212598 443488
rect 4062 443232 4068 443284
rect 4120 443272 4126 443284
rect 213748 443272 213776 443516
rect 215846 443408 215852 443420
rect 4120 443244 213776 443272
rect 214116 443380 215852 443408
rect 4120 443232 4126 443244
rect 3326 443164 3332 443216
rect 3384 443204 3390 443216
rect 214116 443204 214144 443380
rect 215846 443368 215852 443380
rect 215904 443368 215910 443420
rect 3384 443176 214144 443204
rect 216416 443204 216444 443516
rect 220262 443504 220268 443556
rect 220320 443544 220326 443556
rect 224926 443544 224954 443584
rect 220320 443516 224954 443544
rect 220320 443504 220326 443516
rect 234430 443476 234436 443488
rect 224926 443448 234436 443476
rect 216582 443368 216588 443420
rect 216640 443368 216646 443420
rect 217502 443368 217508 443420
rect 217560 443408 217566 443420
rect 224926 443408 224954 443448
rect 234430 443436 234436 443448
rect 234488 443436 234494 443488
rect 234586 443476 234614 443584
rect 239030 443504 239036 443556
rect 239088 443544 239094 443556
rect 240106 443544 240134 443652
rect 242710 443640 242716 443652
rect 242768 443640 242774 443692
rect 248966 443640 248972 443692
rect 249024 443680 249030 443692
rect 297542 443680 297548 443692
rect 249024 443652 297548 443680
rect 249024 443640 249030 443652
rect 297542 443640 297548 443652
rect 297600 443640 297606 443692
rect 239088 443516 240134 443544
rect 241486 443584 259454 443612
rect 239088 443504 239094 443516
rect 241486 443476 241514 443584
rect 242894 443504 242900 443556
rect 242952 443544 242958 443556
rect 242952 443516 256004 443544
rect 242952 443504 242958 443516
rect 234586 443448 241514 443476
rect 242636 443448 245332 443476
rect 217560 443380 224954 443408
rect 217560 443368 217566 443380
rect 225230 443368 225236 443420
rect 225288 443368 225294 443420
rect 225782 443368 225788 443420
rect 225840 443368 225846 443420
rect 226334 443368 226340 443420
rect 226392 443368 226398 443420
rect 228174 443368 228180 443420
rect 228232 443368 228238 443420
rect 229462 443408 229468 443420
rect 229066 443380 229468 443408
rect 216600 443340 216628 443368
rect 225248 443340 225276 443368
rect 216600 443312 225276 443340
rect 220786 443244 222194 443272
rect 220786 443204 220814 443244
rect 216416 443176 220814 443204
rect 222166 443204 222194 443244
rect 225800 443204 225828 443368
rect 222166 443176 225828 443204
rect 3384 443164 3390 443176
rect 3970 443096 3976 443148
rect 4028 443136 4034 443148
rect 226352 443136 226380 443368
rect 4028 443108 226380 443136
rect 4028 443096 4034 443108
rect 4890 443028 4896 443080
rect 4948 443068 4954 443080
rect 228192 443068 228220 443368
rect 4948 443040 212672 443068
rect 4948 443028 4954 443040
rect 3418 442960 3424 443012
rect 3476 443000 3482 443012
rect 212644 443000 212672 443040
rect 212828 443040 228220 443068
rect 212828 443000 212856 443040
rect 229066 443000 229094 443380
rect 229462 443368 229468 443380
rect 229520 443368 229526 443420
rect 233694 443368 233700 443420
rect 233752 443368 233758 443420
rect 239214 443368 239220 443420
rect 239272 443368 239278 443420
rect 239950 443368 239956 443420
rect 240008 443368 240014 443420
rect 3476 442972 212534 443000
rect 212644 442972 212856 443000
rect 212920 442972 229094 443000
rect 233712 443000 233740 443368
rect 239232 443272 239260 443368
rect 239968 443340 239996 443368
rect 239968 443312 240134 443340
rect 240106 443272 240134 443312
rect 242636 443272 242664 443448
rect 242710 443368 242716 443420
rect 242768 443368 242774 443420
rect 239232 443244 239628 443272
rect 240106 443244 242664 443272
rect 239600 443068 239628 443244
rect 242728 443136 242756 443368
rect 245304 443204 245332 443448
rect 254486 443368 254492 443420
rect 254544 443368 254550 443420
rect 254504 443204 254532 443368
rect 245304 443176 254532 443204
rect 255976 443204 256004 443516
rect 256142 443368 256148 443420
rect 256200 443368 256206 443420
rect 259426 443408 259454 443584
rect 265986 443408 265992 443420
rect 259426 443380 265992 443408
rect 265986 443368 265992 443380
rect 266044 443368 266050 443420
rect 256160 443340 256188 443368
rect 298554 443340 298560 443352
rect 256160 443312 298560 443340
rect 298554 443300 298560 443312
rect 298612 443300 298618 443352
rect 266354 443272 266360 443284
rect 259426 443244 266360 443272
rect 259426 443204 259454 443244
rect 266354 443232 266360 443244
rect 266412 443232 266418 443284
rect 255976 443176 259454 443204
rect 265526 443136 265532 443148
rect 242728 443108 265532 443136
rect 265526 443096 265532 443108
rect 265584 443096 265590 443148
rect 266998 443068 267004 443080
rect 239600 443040 267004 443068
rect 266998 443028 267004 443040
rect 267056 443028 267062 443080
rect 298002 443000 298008 443012
rect 233712 442972 298008 443000
rect 3476 442960 3482 442972
rect 212506 442864 212534 442972
rect 212920 442864 212948 442972
rect 298002 442960 298008 442972
rect 298060 442960 298066 443012
rect 212506 442836 212948 442864
rect 266354 440172 266360 440224
rect 266412 440212 266418 440224
rect 298002 440212 298008 440224
rect 266412 440184 298008 440212
rect 266412 440172 266418 440184
rect 298002 440172 298008 440184
rect 298060 440172 298066 440224
rect 265526 436024 265532 436076
rect 265584 436064 265590 436076
rect 297174 436064 297180 436076
rect 265584 436036 297180 436064
rect 265584 436024 265590 436036
rect 297174 436024 297180 436036
rect 297232 436024 297238 436076
rect 267090 431876 267096 431928
rect 267148 431916 267154 431928
rect 298002 431916 298008 431928
rect 267148 431888 298008 431916
rect 267148 431876 267154 431888
rect 298002 431876 298008 431888
rect 298060 431876 298066 431928
rect 384298 431876 384304 431928
rect 384356 431916 384362 431928
rect 580166 431916 580172 431928
rect 384356 431888 580172 431916
rect 384356 431876 384362 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 268470 426368 268476 426420
rect 268528 426408 268534 426420
rect 298002 426408 298008 426420
rect 268528 426380 298008 426408
rect 268528 426368 268534 426380
rect 298002 426368 298008 426380
rect 298060 426368 298066 426420
rect 3142 423580 3148 423632
rect 3200 423620 3206 423632
rect 13078 423620 13084 423632
rect 3200 423592 13084 423620
rect 3200 423580 3206 423592
rect 13078 423580 13084 423592
rect 13136 423580 13142 423632
rect 266998 408416 267004 408468
rect 267056 408456 267062 408468
rect 298002 408456 298008 408468
rect 267056 408428 298008 408456
rect 267056 408416 267062 408428
rect 298002 408416 298008 408428
rect 298060 408416 298066 408468
rect 266170 404268 266176 404320
rect 266228 404308 266234 404320
rect 298002 404308 298008 404320
rect 266228 404280 298008 404308
rect 266228 404268 266234 404280
rect 298002 404268 298008 404280
rect 298060 404268 298066 404320
rect 299566 401208 299572 401260
rect 299624 401248 299630 401260
rect 299624 401220 318794 401248
rect 299624 401208 299630 401220
rect 293862 401072 293868 401124
rect 293920 401112 293926 401124
rect 299658 401112 299664 401124
rect 293920 401084 299664 401112
rect 293920 401072 293926 401084
rect 299658 401072 299664 401084
rect 299716 401072 299722 401124
rect 293770 401004 293776 401056
rect 293828 401044 293834 401056
rect 299474 401044 299480 401056
rect 293828 401016 299480 401044
rect 293828 401004 293834 401016
rect 299474 401004 299480 401016
rect 299532 401004 299538 401056
rect 293586 400936 293592 400988
rect 293644 400976 293650 400988
rect 299566 400976 299572 400988
rect 293644 400948 299572 400976
rect 293644 400936 293650 400948
rect 299566 400936 299572 400948
rect 299624 400936 299630 400988
rect 293678 400868 293684 400920
rect 293736 400908 293742 400920
rect 293736 400880 300256 400908
rect 293736 400868 293742 400880
rect 299566 400732 299572 400784
rect 299624 400772 299630 400784
rect 299842 400772 299848 400784
rect 299624 400744 299848 400772
rect 299624 400732 299630 400744
rect 299842 400732 299848 400744
rect 299900 400732 299906 400784
rect 300228 400772 300256 400880
rect 300228 400744 314654 400772
rect 299474 400664 299480 400716
rect 299532 400704 299538 400716
rect 299532 400676 311940 400704
rect 299532 400664 299538 400676
rect 311912 400648 311940 400676
rect 299658 400596 299664 400648
rect 299716 400636 299722 400648
rect 307570 400636 307576 400648
rect 299716 400608 307576 400636
rect 299716 400596 299722 400608
rect 307570 400596 307576 400608
rect 307628 400596 307634 400648
rect 311894 400596 311900 400648
rect 311952 400596 311958 400648
rect 314626 400636 314654 400744
rect 318766 400704 318794 401220
rect 328426 400880 335354 400908
rect 318766 400676 324268 400704
rect 324240 400648 324268 400676
rect 314626 400608 318794 400636
rect 318766 400568 318794 400608
rect 324222 400596 324228 400648
rect 324280 400596 324286 400648
rect 328426 400568 328454 400880
rect 335326 400636 335354 400880
rect 340966 400636 340972 400648
rect 335326 400608 340972 400636
rect 340966 400596 340972 400608
rect 341024 400596 341030 400648
rect 318766 400540 328454 400568
rect 298554 400120 298560 400172
rect 298612 400160 298618 400172
rect 579982 400160 579988 400172
rect 298612 400132 579988 400160
rect 298612 400120 298618 400132
rect 579982 400120 579988 400132
rect 580040 400120 580046 400172
rect 293310 400052 293316 400104
rect 293368 400092 293374 400104
rect 385034 400092 385040 400104
rect 293368 400064 385040 400092
rect 293368 400052 293374 400064
rect 385034 400052 385040 400064
rect 385092 400052 385098 400104
rect 217226 399168 217232 399220
rect 217284 399208 217290 399220
rect 217284 399180 217364 399208
rect 217284 399168 217290 399180
rect 216950 399032 216956 399084
rect 217008 399072 217014 399084
rect 217226 399072 217232 399084
rect 217008 399044 217232 399072
rect 217008 399032 217014 399044
rect 217226 399032 217232 399044
rect 217284 399032 217290 399084
rect 217336 398868 217364 399180
rect 244366 399100 244372 399152
rect 244424 399140 244430 399152
rect 437474 399140 437480 399152
rect 244424 399112 437480 399140
rect 244424 399100 244430 399112
rect 437474 399100 437480 399112
rect 437532 399100 437538 399152
rect 238726 399044 253612 399072
rect 217594 398964 217600 399016
rect 217652 399004 217658 399016
rect 217652 398976 217824 399004
rect 217652 398964 217658 398976
rect 217686 398936 217692 398948
rect 217152 398840 217364 398868
rect 217520 398908 217692 398936
rect 208026 398760 208032 398812
rect 208084 398800 208090 398812
rect 210050 398800 210056 398812
rect 208084 398772 210056 398800
rect 208084 398760 208090 398772
rect 210050 398760 210056 398772
rect 210108 398760 210114 398812
rect 210234 398760 210240 398812
rect 210292 398800 210298 398812
rect 210292 398772 214696 398800
rect 210292 398760 210298 398772
rect 207658 398692 207664 398744
rect 207716 398732 207722 398744
rect 207716 398704 214604 398732
rect 207716 398692 207722 398704
rect 207934 398624 207940 398676
rect 207992 398664 207998 398676
rect 210142 398664 210148 398676
rect 207992 398636 210148 398664
rect 207992 398624 207998 398636
rect 210142 398624 210148 398636
rect 210200 398624 210206 398676
rect 214006 398624 214012 398676
rect 214064 398664 214070 398676
rect 214466 398664 214472 398676
rect 214064 398636 214472 398664
rect 214064 398624 214070 398636
rect 214466 398624 214472 398636
rect 214524 398624 214530 398676
rect 207014 398556 207020 398608
rect 207072 398596 207078 398608
rect 207072 398568 214512 398596
rect 207072 398556 207078 398568
rect 207842 398488 207848 398540
rect 207900 398528 207906 398540
rect 210234 398528 210240 398540
rect 207900 398500 210240 398528
rect 207900 398488 207906 398500
rect 210234 398488 210240 398500
rect 210292 398488 210298 398540
rect 203518 398420 203524 398472
rect 203576 398460 203582 398472
rect 211798 398460 211804 398472
rect 203576 398432 211804 398460
rect 203576 398420 203582 398432
rect 211798 398420 211804 398432
rect 211856 398420 211862 398472
rect 209222 398352 209228 398404
rect 209280 398392 209286 398404
rect 212166 398392 212172 398404
rect 209280 398364 212172 398392
rect 209280 398352 209286 398364
rect 212166 398352 212172 398364
rect 212224 398352 212230 398404
rect 214484 398392 214512 398568
rect 214576 398460 214604 398704
rect 214668 398664 214696 398772
rect 217152 398664 217180 398840
rect 217520 398744 217548 398908
rect 217686 398896 217692 398908
rect 217744 398896 217750 398948
rect 217502 398692 217508 398744
rect 217560 398692 217566 398744
rect 217594 398692 217600 398744
rect 217652 398732 217658 398744
rect 217796 398732 217824 398976
rect 219342 398964 219348 399016
rect 219400 399004 219406 399016
rect 219434 399004 219440 399016
rect 219400 398976 219440 399004
rect 219400 398964 219406 398976
rect 219434 398964 219440 398976
rect 219492 398964 219498 399016
rect 236086 398896 236092 398948
rect 236144 398936 236150 398948
rect 238726 398936 238754 399044
rect 253584 398936 253612 399044
rect 253658 399032 253664 399084
rect 253716 399072 253722 399084
rect 277394 399072 277400 399084
rect 253716 399044 277400 399072
rect 253716 399032 253722 399044
rect 277394 399032 277400 399044
rect 277452 399032 277458 399084
rect 256050 398964 256056 399016
rect 256108 399004 256114 399016
rect 299474 399004 299480 399016
rect 256108 398976 299480 399004
rect 256108 398964 256114 398976
rect 299474 398964 299480 398976
rect 299532 398964 299538 399016
rect 331214 398936 331220 398948
rect 236144 398908 238754 398936
rect 241486 398908 251174 398936
rect 253584 398908 331220 398936
rect 236144 398896 236150 398908
rect 230842 398760 230848 398812
rect 230900 398800 230906 398812
rect 241486 398800 241514 398908
rect 251146 398868 251174 398908
rect 331214 398896 331220 398908
rect 331272 398896 331278 398948
rect 263594 398868 263600 398880
rect 230900 398772 241514 398800
rect 244752 398840 248092 398868
rect 251146 398840 263600 398868
rect 230900 398760 230906 398772
rect 217652 398704 217824 398732
rect 217652 398692 217658 398704
rect 217226 398664 217232 398676
rect 214668 398636 215294 398664
rect 217152 398636 217232 398664
rect 215266 398528 215294 398636
rect 217226 398624 217232 398636
rect 217284 398624 217290 398676
rect 217778 398664 217784 398676
rect 217336 398636 217784 398664
rect 217336 398528 217364 398636
rect 217778 398624 217784 398636
rect 217836 398624 217842 398676
rect 229278 398624 229284 398676
rect 229336 398664 229342 398676
rect 230014 398664 230020 398676
rect 229336 398636 230020 398664
rect 229336 398624 229342 398636
rect 230014 398624 230020 398636
rect 230072 398624 230078 398676
rect 244752 398664 244780 398840
rect 244826 398692 244832 398744
rect 244884 398732 244890 398744
rect 248064 398732 248092 398840
rect 263594 398828 263600 398840
rect 263652 398828 263658 398880
rect 296622 398760 296628 398812
rect 296680 398800 296686 398812
rect 379238 398800 379244 398812
rect 296680 398772 379244 398800
rect 296680 398760 296686 398772
rect 379238 398760 379244 398772
rect 379296 398760 379302 398812
rect 256050 398732 256056 398744
rect 244884 398704 247816 398732
rect 248064 398704 256056 398732
rect 244884 398692 244890 398704
rect 238726 398636 244780 398664
rect 215266 398500 217364 398528
rect 217778 398488 217784 398540
rect 217836 398528 217842 398540
rect 222838 398528 222844 398540
rect 217836 398500 222844 398528
rect 217836 398488 217842 398500
rect 222838 398488 222844 398500
rect 222896 398488 222902 398540
rect 228450 398488 228456 398540
rect 228508 398528 228514 398540
rect 230014 398528 230020 398540
rect 228508 398500 230020 398528
rect 228508 398488 228514 398500
rect 230014 398488 230020 398500
rect 230072 398488 230078 398540
rect 233602 398488 233608 398540
rect 233660 398528 233666 398540
rect 238726 398528 238754 398636
rect 239858 398556 239864 398608
rect 239916 398596 239922 398608
rect 245654 398596 245660 398608
rect 239916 398568 245660 398596
rect 239916 398556 239922 398568
rect 245654 398556 245660 398568
rect 245712 398556 245718 398608
rect 247788 398596 247816 398704
rect 256050 398692 256056 398704
rect 256108 398692 256114 398744
rect 295886 398692 295892 398744
rect 295944 398732 295950 398744
rect 303890 398732 303896 398744
rect 295944 398704 303896 398732
rect 295944 398692 295950 398704
rect 303890 398692 303896 398704
rect 303948 398692 303954 398744
rect 255498 398624 255504 398676
rect 255556 398664 255562 398676
rect 269758 398664 269764 398676
rect 255556 398636 269764 398664
rect 255556 398624 255562 398636
rect 269758 398624 269764 398636
rect 269816 398624 269822 398676
rect 299566 398624 299572 398676
rect 299624 398664 299630 398676
rect 374730 398664 374736 398676
rect 299624 398636 374736 398664
rect 299624 398624 299630 398636
rect 374730 398624 374736 398636
rect 374788 398624 374794 398676
rect 261478 398596 261484 398608
rect 247788 398568 261484 398596
rect 261478 398556 261484 398568
rect 261536 398556 261542 398608
rect 293218 398556 293224 398608
rect 293276 398596 293282 398608
rect 366358 398596 366364 398608
rect 293276 398568 366364 398596
rect 293276 398556 293282 398568
rect 366358 398556 366364 398568
rect 366416 398556 366422 398608
rect 233660 398500 238754 398528
rect 233660 398488 233666 398500
rect 245930 398488 245936 398540
rect 245988 398528 245994 398540
rect 264238 398528 264244 398540
rect 245988 398500 264244 398528
rect 245988 398488 245994 398500
rect 264238 398488 264244 398500
rect 264296 398488 264302 398540
rect 299382 398488 299388 398540
rect 299440 398528 299446 398540
rect 370866 398528 370872 398540
rect 299440 398500 370872 398528
rect 299440 398488 299446 398500
rect 370866 398488 370872 398500
rect 370924 398488 370930 398540
rect 223390 398460 223396 398472
rect 214576 398432 223396 398460
rect 223390 398420 223396 398432
rect 223448 398420 223454 398472
rect 233326 398420 233332 398472
rect 233384 398460 233390 398472
rect 239858 398460 239864 398472
rect 233384 398432 239864 398460
rect 233384 398420 233390 398432
rect 239858 398420 239864 398432
rect 239916 398420 239922 398472
rect 240410 398420 240416 398472
rect 240468 398460 240474 398472
rect 245378 398460 245384 398472
rect 240468 398432 245384 398460
rect 240468 398420 240474 398432
rect 245378 398420 245384 398432
rect 245436 398420 245442 398472
rect 246206 398420 246212 398472
rect 246264 398460 246270 398472
rect 264330 398460 264336 398472
rect 246264 398432 264336 398460
rect 246264 398420 246270 398432
rect 264330 398420 264336 398432
rect 264388 398420 264394 398472
rect 296530 398420 296536 398472
rect 296588 398460 296594 398472
rect 362494 398460 362500 398472
rect 296588 398432 362500 398460
rect 296588 398420 296594 398432
rect 362494 398420 362500 398432
rect 362552 398420 362558 398472
rect 226426 398392 226432 398404
rect 214484 398364 226432 398392
rect 226426 398352 226432 398364
rect 226484 398352 226490 398404
rect 238726 398364 255360 398392
rect 204898 398284 204904 398336
rect 204956 398324 204962 398336
rect 212258 398324 212264 398336
rect 204956 398296 212264 398324
rect 204956 398284 204962 398296
rect 212258 398284 212264 398296
rect 212316 398284 212322 398336
rect 213362 398284 213368 398336
rect 213420 398324 213426 398336
rect 223114 398324 223120 398336
rect 213420 398296 223120 398324
rect 213420 398284 213426 398296
rect 223114 398284 223120 398296
rect 223172 398284 223178 398336
rect 229738 398284 229744 398336
rect 229796 398324 229802 398336
rect 238726 398324 238754 398364
rect 229796 398296 238754 398324
rect 229796 398284 229802 398296
rect 241514 398284 241520 398336
rect 241572 398324 241578 398336
rect 249058 398324 249064 398336
rect 241572 398296 249064 398324
rect 241572 398284 241578 398296
rect 249058 398284 249064 398296
rect 249116 398284 249122 398336
rect 252646 398284 252652 398336
rect 252704 398324 252710 398336
rect 252704 398296 255268 398324
rect 252704 398284 252710 398296
rect 171134 398216 171140 398268
rect 171192 398256 171198 398268
rect 223666 398256 223672 398268
rect 171192 398228 223672 398256
rect 171192 398216 171198 398228
rect 223666 398216 223672 398228
rect 223724 398216 223730 398268
rect 230566 398216 230572 398268
rect 230624 398256 230630 398268
rect 230624 398228 253934 398256
rect 230624 398216 230630 398228
rect 125594 398148 125600 398200
rect 125652 398188 125658 398200
rect 220078 398188 220084 398200
rect 125652 398160 220084 398188
rect 125652 398148 125658 398160
rect 220078 398148 220084 398160
rect 220136 398148 220142 398200
rect 242066 398148 242072 398200
rect 242124 398188 242130 398200
rect 242124 398160 244228 398188
rect 242124 398148 242130 398160
rect 24854 398080 24860 398132
rect 24912 398120 24918 398132
rect 204898 398120 204904 398132
rect 24912 398092 204904 398120
rect 24912 398080 24918 398092
rect 204898 398080 204904 398092
rect 204956 398080 204962 398132
rect 209774 398080 209780 398132
rect 209832 398120 209838 398132
rect 210694 398120 210700 398132
rect 209832 398092 210700 398120
rect 209832 398080 209838 398092
rect 210694 398080 210700 398092
rect 210752 398080 210758 398132
rect 212442 398080 212448 398132
rect 212500 398120 212506 398132
rect 225046 398120 225052 398132
rect 212500 398092 225052 398120
rect 212500 398080 212506 398092
rect 225046 398080 225052 398092
rect 225104 398080 225110 398132
rect 210142 398012 210148 398064
rect 210200 398052 210206 398064
rect 218330 398052 218336 398064
rect 210200 398024 218336 398052
rect 210200 398012 210206 398024
rect 218330 398012 218336 398024
rect 218388 398012 218394 398064
rect 210050 397944 210056 397996
rect 210108 397984 210114 397996
rect 218882 397984 218888 397996
rect 210108 397956 218888 397984
rect 210108 397944 210114 397956
rect 218882 397944 218888 397956
rect 218940 397944 218946 397996
rect 238202 397944 238208 397996
rect 238260 397984 238266 397996
rect 238260 397956 238754 397984
rect 238260 397944 238266 397956
rect 211522 397876 211528 397928
rect 211580 397916 211586 397928
rect 217226 397916 217232 397928
rect 211580 397888 217232 397916
rect 211580 397876 211586 397888
rect 217226 397876 217232 397888
rect 217284 397876 217290 397928
rect 219434 397876 219440 397928
rect 219492 397876 219498 397928
rect 238726 397916 238754 397956
rect 239306 397944 239312 397996
rect 239364 397984 239370 397996
rect 242618 397984 242624 397996
rect 239364 397956 242624 397984
rect 239364 397944 239370 397956
rect 242618 397944 242624 397956
rect 242676 397944 242682 397996
rect 244200 397984 244228 398160
rect 245654 398080 245660 398132
rect 245712 398120 245718 398132
rect 246482 398120 246488 398132
rect 245712 398092 246488 398120
rect 245712 398080 245718 398092
rect 246482 398080 246488 398092
rect 246540 398080 246546 398132
rect 247678 398080 247684 398132
rect 247736 398120 247742 398132
rect 247954 398120 247960 398132
rect 247736 398092 247960 398120
rect 247736 398080 247742 398092
rect 247954 398080 247960 398092
rect 248012 398080 248018 398132
rect 244274 398012 244280 398064
rect 244332 398052 244338 398064
rect 253906 398052 253934 398228
rect 255240 398188 255268 398296
rect 255332 398256 255360 398364
rect 255590 398352 255596 398404
rect 255648 398392 255654 398404
rect 275370 398392 275376 398404
rect 255648 398364 275376 398392
rect 255648 398352 255654 398364
rect 275370 398352 275376 398364
rect 275428 398352 275434 398404
rect 295794 398352 295800 398404
rect 295852 398392 295858 398404
rect 357986 398392 357992 398404
rect 295852 398364 357992 398392
rect 295852 398352 295858 398364
rect 357986 398352 357992 398364
rect 358044 398352 358050 398404
rect 257522 398284 257528 398336
rect 257580 398324 257586 398336
rect 264974 398324 264980 398336
rect 257580 398296 264980 398324
rect 257580 398284 257586 398296
rect 264974 398284 264980 398296
rect 265032 398284 265038 398336
rect 293494 398284 293500 398336
rect 293552 398324 293558 398336
rect 349614 398324 349620 398336
rect 293552 398296 349620 398324
rect 293552 398284 293558 398296
rect 349614 398284 349620 398296
rect 349672 398284 349678 398336
rect 256694 398256 256700 398268
rect 255332 398228 256700 398256
rect 256694 398216 256700 398228
rect 256752 398216 256758 398268
rect 298646 398216 298652 398268
rect 298704 398256 298710 398268
rect 329006 398256 329012 398268
rect 298704 398228 329012 398256
rect 298704 398216 298710 398228
rect 329006 398216 329012 398228
rect 329064 398216 329070 398268
rect 543734 398188 543740 398200
rect 255240 398160 543740 398188
rect 543734 398148 543740 398160
rect 543792 398148 543798 398200
rect 254302 398080 254308 398132
rect 254360 398120 254366 398132
rect 564434 398120 564440 398132
rect 254360 398092 564440 398120
rect 254360 398080 254366 398092
rect 564434 398080 564440 398092
rect 564492 398080 564498 398132
rect 259546 398052 259552 398064
rect 244332 398024 249196 398052
rect 253906 398024 259552 398052
rect 244332 398012 244338 398024
rect 249168 397984 249196 398024
rect 259546 398012 259552 398024
rect 259604 398012 259610 398064
rect 293402 398012 293408 398064
rect 293460 398052 293466 398064
rect 320634 398052 320640 398064
rect 293460 398024 320640 398052
rect 293460 398012 293466 398024
rect 320634 398012 320640 398024
rect 320692 398012 320698 398064
rect 258810 397984 258816 397996
rect 244200 397956 249104 397984
rect 249168 397956 258816 397984
rect 238726 397888 239444 397916
rect 206278 397808 206284 397860
rect 206336 397848 206342 397860
rect 219452 397848 219480 397876
rect 206336 397820 219480 397848
rect 206336 397808 206342 397820
rect 236362 397808 236368 397860
rect 236420 397848 236426 397860
rect 239306 397848 239312 397860
rect 236420 397820 239312 397848
rect 236420 397808 236426 397820
rect 239306 397808 239312 397820
rect 239364 397808 239370 397860
rect 210234 397740 210240 397792
rect 210292 397780 210298 397792
rect 216950 397780 216956 397792
rect 210292 397752 216956 397780
rect 210292 397740 210298 397752
rect 216950 397740 216956 397752
rect 217008 397740 217014 397792
rect 217042 397740 217048 397792
rect 217100 397780 217106 397792
rect 217778 397780 217784 397792
rect 217100 397752 217784 397780
rect 217100 397740 217106 397752
rect 217778 397740 217784 397752
rect 217836 397740 217842 397792
rect 219434 397740 219440 397792
rect 219492 397780 219498 397792
rect 227438 397780 227444 397792
rect 219492 397752 227444 397780
rect 219492 397740 219498 397752
rect 227438 397740 227444 397752
rect 227496 397740 227502 397792
rect 193214 397672 193220 397724
rect 193272 397712 193278 397724
rect 225322 397712 225328 397724
rect 193272 397684 200114 397712
rect 193272 397672 193278 397684
rect 200086 397644 200114 397684
rect 210896 397684 225328 397712
rect 210896 397644 210924 397684
rect 225322 397672 225328 397684
rect 225380 397672 225386 397724
rect 228266 397672 228272 397724
rect 228324 397712 228330 397724
rect 230474 397712 230480 397724
rect 228324 397684 230480 397712
rect 228324 397672 228330 397684
rect 230474 397672 230480 397684
rect 230532 397672 230538 397724
rect 231946 397672 231952 397724
rect 232004 397712 232010 397724
rect 239416 397712 239444 397888
rect 244826 397876 244832 397928
rect 244884 397916 244890 397928
rect 245930 397916 245936 397928
rect 244884 397888 245936 397916
rect 244884 397876 244890 397888
rect 245930 397876 245936 397888
rect 245988 397876 245994 397928
rect 243170 397808 243176 397860
rect 243228 397848 243234 397860
rect 249076 397848 249104 397956
rect 258810 397944 258816 397956
rect 258868 397944 258874 397996
rect 266078 397944 266084 397996
rect 266136 397984 266142 397996
rect 316126 397984 316132 397996
rect 266136 397956 316132 397984
rect 266136 397944 266142 397956
rect 316126 397944 316132 397956
rect 316184 397944 316190 397996
rect 264974 397876 264980 397928
rect 265032 397916 265038 397928
rect 345750 397916 345756 397928
rect 265032 397888 345756 397916
rect 265032 397876 265038 397888
rect 345750 397876 345756 397888
rect 345808 397876 345814 397928
rect 256418 397848 256424 397860
rect 243228 397820 249012 397848
rect 249076 397820 256424 397848
rect 243228 397808 243234 397820
rect 243722 397740 243728 397792
rect 243780 397780 243786 397792
rect 248984 397780 249012 397820
rect 256418 397808 256424 397820
rect 256476 397808 256482 397860
rect 256602 397780 256608 397792
rect 243780 397752 245700 397780
rect 248984 397752 256608 397780
rect 243780 397740 243786 397752
rect 244826 397712 244832 397724
rect 232004 397684 238754 397712
rect 239416 397684 244832 397712
rect 232004 397672 232010 397684
rect 200086 397616 210924 397644
rect 217778 397604 217784 397656
rect 217836 397644 217842 397656
rect 220814 397644 220820 397656
rect 217836 397616 220820 397644
rect 217836 397604 217842 397616
rect 220814 397604 220820 397616
rect 220872 397604 220878 397656
rect 222194 397604 222200 397656
rect 222252 397644 222258 397656
rect 227622 397644 227628 397656
rect 222252 397616 227628 397644
rect 222252 397604 222258 397616
rect 227622 397604 227628 397616
rect 227680 397604 227686 397656
rect 234062 397604 234068 397656
rect 234120 397604 234126 397656
rect 238726 397644 238754 397684
rect 244826 397672 244832 397684
rect 244884 397672 244890 397724
rect 244458 397644 244464 397656
rect 238726 397616 244464 397644
rect 244458 397604 244464 397616
rect 244516 397604 244522 397656
rect 245672 397644 245700 397752
rect 256602 397740 256608 397752
rect 256660 397740 256666 397792
rect 245930 397672 245936 397724
rect 245988 397712 245994 397724
rect 246758 397712 246764 397724
rect 245988 397684 246764 397712
rect 245988 397672 245994 397684
rect 246758 397672 246764 397684
rect 246816 397672 246822 397724
rect 249058 397672 249064 397724
rect 249116 397712 249122 397724
rect 256510 397712 256516 397724
rect 249116 397684 256516 397712
rect 249116 397672 249122 397684
rect 256510 397672 256516 397684
rect 256568 397672 256574 397724
rect 257614 397644 257620 397656
rect 245672 397616 257620 397644
rect 257614 397604 257620 397616
rect 257672 397604 257678 397656
rect 209038 397536 209044 397588
rect 209096 397576 209102 397588
rect 210786 397576 210792 397588
rect 209096 397548 210792 397576
rect 209096 397536 209102 397548
rect 210786 397536 210792 397548
rect 210844 397536 210850 397588
rect 211522 397576 211528 397588
rect 210896 397548 211528 397576
rect 210234 397468 210240 397520
rect 210292 397508 210298 397520
rect 210694 397508 210700 397520
rect 210292 397480 210700 397508
rect 210292 397468 210298 397480
rect 210694 397468 210700 397480
rect 210752 397468 210758 397520
rect 210896 397508 210924 397548
rect 211522 397536 211528 397548
rect 211580 397536 211586 397588
rect 211890 397536 211896 397588
rect 211948 397576 211954 397588
rect 215018 397576 215024 397588
rect 211948 397548 215024 397576
rect 211948 397536 211954 397548
rect 215018 397536 215024 397548
rect 215076 397536 215082 397588
rect 218790 397576 218796 397588
rect 215128 397548 218796 397576
rect 210804 397480 210924 397508
rect 210804 397452 210832 397480
rect 211154 397468 211160 397520
rect 211212 397508 211218 397520
rect 213546 397508 213552 397520
rect 211212 397480 213552 397508
rect 211212 397468 211218 397480
rect 213546 397468 213552 397480
rect 213604 397468 213610 397520
rect 210786 397400 210792 397452
rect 210844 397400 210850 397452
rect 215018 397400 215024 397452
rect 215076 397440 215082 397452
rect 215128 397440 215156 397548
rect 218790 397536 218796 397548
rect 218848 397536 218854 397588
rect 218882 397536 218888 397588
rect 218940 397576 218946 397588
rect 220722 397576 220728 397588
rect 218940 397548 220728 397576
rect 218940 397536 218946 397548
rect 220722 397536 220728 397548
rect 220780 397536 220786 397588
rect 224954 397536 224960 397588
rect 225012 397576 225018 397588
rect 227162 397576 227168 397588
rect 225012 397548 227168 397576
rect 225012 397536 225018 397548
rect 227162 397536 227168 397548
rect 227220 397536 227226 397588
rect 234080 397576 234108 397604
rect 234080 397548 234384 397576
rect 234356 397520 234384 397548
rect 239306 397536 239312 397588
rect 239364 397576 239370 397588
rect 240042 397576 240048 397588
rect 239364 397548 240048 397576
rect 239364 397536 239370 397548
rect 240042 397536 240048 397548
rect 240100 397536 240106 397588
rect 240888 397548 242756 397576
rect 220078 397468 220084 397520
rect 220136 397508 220142 397520
rect 222378 397508 222384 397520
rect 220136 397480 222384 397508
rect 220136 397468 220142 397480
rect 222378 397468 222384 397480
rect 222436 397468 222442 397520
rect 225046 397468 225052 397520
rect 225104 397508 225110 397520
rect 225598 397508 225604 397520
rect 225104 397480 225604 397508
rect 225104 397468 225110 397480
rect 225598 397468 225604 397480
rect 225656 397468 225662 397520
rect 226426 397468 226432 397520
rect 226484 397508 226490 397520
rect 227714 397508 227720 397520
rect 226484 397480 227720 397508
rect 226484 397468 226490 397480
rect 227714 397468 227720 397480
rect 227772 397468 227778 397520
rect 231486 397468 231492 397520
rect 231544 397508 231550 397520
rect 234062 397508 234068 397520
rect 231544 397480 234068 397508
rect 231544 397468 231550 397480
rect 234062 397468 234068 397480
rect 234120 397468 234126 397520
rect 234338 397468 234344 397520
rect 234396 397468 234402 397520
rect 238754 397468 238760 397520
rect 238812 397508 238818 397520
rect 240888 397508 240916 397548
rect 238812 397480 240916 397508
rect 238812 397468 238818 397480
rect 240962 397468 240968 397520
rect 241020 397508 241026 397520
rect 242618 397508 242624 397520
rect 241020 397480 242624 397508
rect 241020 397468 241026 397480
rect 242618 397468 242624 397480
rect 242676 397468 242682 397520
rect 242728 397508 242756 397548
rect 248782 397536 248788 397588
rect 248840 397576 248846 397588
rect 257430 397576 257436 397588
rect 248840 397548 253796 397576
rect 248840 397536 248846 397548
rect 243998 397508 244004 397520
rect 242728 397480 244004 397508
rect 243998 397468 244004 397480
rect 244056 397468 244062 397520
rect 244458 397468 244464 397520
rect 244516 397508 244522 397520
rect 253658 397508 253664 397520
rect 244516 397480 253664 397508
rect 244516 397468 244522 397480
rect 253658 397468 253664 397480
rect 253716 397468 253722 397520
rect 253768 397508 253796 397548
rect 253952 397548 257436 397576
rect 253768 397480 253888 397508
rect 215076 397412 215156 397440
rect 215076 397400 215082 397412
rect 217226 397400 217232 397452
rect 217284 397440 217290 397452
rect 226610 397440 226616 397452
rect 217284 397412 226616 397440
rect 217284 397400 217290 397412
rect 226610 397400 226616 397412
rect 226668 397400 226674 397452
rect 253860 397440 253888 397480
rect 253952 397440 253980 397548
rect 257430 397536 257436 397548
rect 257488 397536 257494 397588
rect 254026 397468 254032 397520
rect 254084 397508 254090 397520
rect 256326 397508 256332 397520
rect 254084 397480 256332 397508
rect 254084 397468 254090 397480
rect 256326 397468 256332 397480
rect 256384 397468 256390 397520
rect 253860 397412 253980 397440
rect 211614 397332 211620 397384
rect 211672 397372 211678 397384
rect 218606 397372 218612 397384
rect 211672 397344 218612 397372
rect 211672 397332 211678 397344
rect 218606 397332 218612 397344
rect 218664 397332 218670 397384
rect 226058 397372 226064 397384
rect 218716 397344 226064 397372
rect 201494 397264 201500 397316
rect 201552 397304 201558 397316
rect 218716 397304 218744 397344
rect 226058 397332 226064 397344
rect 226116 397332 226122 397384
rect 225506 397304 225512 397316
rect 201552 397276 218744 397304
rect 224926 397276 225512 397304
rect 201552 397264 201558 397276
rect 212534 397196 212540 397248
rect 212592 397236 212598 397248
rect 213454 397236 213460 397248
rect 212592 397208 213460 397236
rect 212592 397196 212598 397208
rect 213454 397196 213460 397208
rect 213512 397196 213518 397248
rect 194594 397128 194600 397180
rect 194652 397168 194658 397180
rect 224926 397168 224954 397276
rect 225506 397264 225512 397276
rect 225564 397264 225570 397316
rect 247034 397196 247040 397248
rect 247092 397236 247098 397248
rect 247586 397236 247592 397248
rect 247092 397208 247592 397236
rect 247092 397196 247098 397208
rect 247586 397196 247592 397208
rect 247644 397196 247650 397248
rect 247678 397196 247684 397248
rect 247736 397236 247742 397248
rect 256142 397236 256148 397248
rect 247736 397208 256148 397236
rect 247736 397196 247742 397208
rect 256142 397196 256148 397208
rect 256200 397196 256206 397248
rect 194652 397140 224954 397168
rect 194652 397128 194658 397140
rect 227806 397128 227812 397180
rect 227864 397168 227870 397180
rect 229002 397168 229008 397180
rect 227864 397140 229008 397168
rect 227864 397128 227870 397140
rect 229002 397128 229008 397140
rect 229060 397128 229066 397180
rect 235442 397128 235448 397180
rect 235500 397168 235506 397180
rect 235626 397168 235632 397180
rect 235500 397140 235632 397168
rect 235500 397128 235506 397140
rect 235626 397128 235632 397140
rect 235684 397128 235690 397180
rect 238754 397128 238760 397180
rect 238812 397168 238818 397180
rect 239398 397168 239404 397180
rect 238812 397140 239404 397168
rect 238812 397128 238818 397140
rect 239398 397128 239404 397140
rect 239456 397128 239462 397180
rect 241698 397128 241704 397180
rect 241756 397168 241762 397180
rect 249058 397168 249064 397180
rect 241756 397140 249064 397168
rect 241756 397128 241762 397140
rect 249058 397128 249064 397140
rect 249116 397128 249122 397180
rect 256050 397168 256056 397180
rect 249720 397140 256056 397168
rect 160094 397060 160100 397112
rect 160152 397100 160158 397112
rect 222746 397100 222752 397112
rect 160152 397072 222752 397100
rect 160152 397060 160158 397072
rect 222746 397060 222752 397072
rect 222804 397060 222810 397112
rect 246206 397060 246212 397112
rect 246264 397100 246270 397112
rect 249720 397100 249748 397140
rect 256050 397128 256056 397140
rect 256108 397128 256114 397180
rect 246264 397072 249748 397100
rect 246264 397060 246270 397072
rect 144914 396992 144920 397044
rect 144972 397032 144978 397044
rect 221642 397032 221648 397044
rect 144972 397004 221648 397032
rect 144972 396992 144978 397004
rect 221642 396992 221648 397004
rect 221700 396992 221706 397044
rect 227806 396992 227812 397044
rect 227864 397032 227870 397044
rect 228726 397032 228732 397044
rect 227864 397004 228732 397032
rect 227864 396992 227870 397004
rect 228726 396992 228732 397004
rect 228784 396992 228790 397044
rect 231854 396992 231860 397044
rect 231912 397032 231918 397044
rect 232866 397032 232872 397044
rect 231912 397004 232872 397032
rect 231912 396992 231918 397004
rect 232866 396992 232872 397004
rect 232924 396992 232930 397044
rect 234890 396992 234896 397044
rect 234948 397032 234954 397044
rect 235442 397032 235448 397044
rect 234948 397004 235448 397032
rect 234948 396992 234954 397004
rect 235442 396992 235448 397004
rect 235500 396992 235506 397044
rect 238846 396992 238852 397044
rect 238904 397032 238910 397044
rect 239398 397032 239404 397044
rect 238904 397004 239404 397032
rect 238904 396992 238910 397004
rect 239398 396992 239404 397004
rect 239456 396992 239462 397044
rect 242176 397004 244780 397032
rect 135254 396924 135260 396976
rect 135312 396964 135318 396976
rect 217778 396964 217784 396976
rect 135312 396936 217784 396964
rect 135312 396924 135318 396936
rect 217778 396924 217784 396936
rect 217836 396924 217842 396976
rect 229738 396924 229744 396976
rect 229796 396964 229802 396976
rect 229796 396936 234108 396964
rect 229796 396924 229802 396936
rect 131114 396856 131120 396908
rect 131172 396896 131178 396908
rect 220538 396896 220544 396908
rect 131172 396868 220544 396896
rect 131172 396856 131178 396868
rect 220538 396856 220544 396868
rect 220596 396856 220602 396908
rect 228082 396856 228088 396908
rect 228140 396896 228146 396908
rect 228726 396896 228732 396908
rect 228140 396868 228732 396896
rect 228140 396856 228146 396868
rect 228726 396856 228732 396868
rect 228784 396856 228790 396908
rect 230566 396856 230572 396908
rect 230624 396896 230630 396908
rect 231578 396896 231584 396908
rect 230624 396868 231584 396896
rect 230624 396856 230630 396868
rect 231578 396856 231584 396868
rect 231636 396856 231642 396908
rect 231854 396856 231860 396908
rect 231912 396896 231918 396908
rect 232498 396896 232504 396908
rect 231912 396868 232504 396896
rect 231912 396856 231918 396868
rect 232498 396856 232504 396868
rect 232556 396856 232562 396908
rect 233326 396856 233332 396908
rect 233384 396896 233390 396908
rect 233694 396896 233700 396908
rect 233384 396868 233700 396896
rect 233384 396856 233390 396868
rect 233694 396856 233700 396868
rect 233752 396856 233758 396908
rect 106274 396788 106280 396840
rect 106332 396828 106338 396840
rect 211614 396828 211620 396840
rect 106332 396800 211620 396828
rect 106332 396788 106338 396800
rect 211614 396788 211620 396800
rect 211672 396788 211678 396840
rect 212718 396788 212724 396840
rect 212776 396828 212782 396840
rect 213178 396828 213184 396840
rect 212776 396800 213184 396828
rect 212776 396788 212782 396800
rect 213178 396788 213184 396800
rect 213236 396788 213242 396840
rect 229370 396788 229376 396840
rect 229428 396828 229434 396840
rect 230106 396828 230112 396840
rect 229428 396800 230112 396828
rect 229428 396788 229434 396800
rect 230106 396788 230112 396800
rect 230164 396788 230170 396840
rect 231946 396788 231952 396840
rect 232004 396828 232010 396840
rect 232314 396828 232320 396840
rect 232004 396800 232320 396828
rect 232004 396788 232010 396800
rect 232314 396788 232320 396800
rect 232372 396788 232378 396840
rect 234080 396828 234108 396936
rect 237374 396924 237380 396976
rect 237432 396964 237438 396976
rect 238386 396964 238392 396976
rect 237432 396936 238392 396964
rect 237432 396924 237438 396936
rect 238386 396924 238392 396936
rect 238444 396924 238450 396976
rect 238938 396924 238944 396976
rect 238996 396964 239002 396976
rect 239306 396964 239312 396976
rect 238996 396936 239312 396964
rect 238996 396924 239002 396936
rect 239306 396924 239312 396936
rect 239364 396924 239370 396976
rect 240778 396924 240784 396976
rect 240836 396964 240842 396976
rect 241422 396964 241428 396976
rect 240836 396936 241428 396964
rect 240836 396924 240842 396936
rect 241422 396924 241428 396936
rect 241480 396924 241486 396976
rect 234614 396856 234620 396908
rect 234672 396896 234678 396908
rect 234982 396896 234988 396908
rect 234672 396868 234988 396896
rect 234672 396856 234678 396868
rect 234982 396856 234988 396868
rect 235040 396856 235046 396908
rect 237006 396856 237012 396908
rect 237064 396896 237070 396908
rect 242176 396896 242204 397004
rect 237064 396868 242204 396896
rect 237064 396856 237070 396868
rect 242250 396856 242256 396908
rect 242308 396896 242314 396908
rect 244752 396896 244780 397004
rect 342254 396896 342260 396908
rect 242308 396868 244228 396896
rect 244752 396868 342260 396896
rect 242308 396856 242314 396868
rect 242434 396828 242440 396840
rect 234080 396800 242440 396828
rect 242434 396788 242440 396800
rect 242492 396788 242498 396840
rect 242802 396788 242808 396840
rect 242860 396828 242866 396840
rect 243538 396828 243544 396840
rect 242860 396800 243544 396828
rect 242860 396788 242866 396800
rect 243538 396788 243544 396800
rect 243596 396788 243602 396840
rect 244200 396828 244228 396868
rect 342254 396856 342260 396868
rect 342312 396856 342318 396908
rect 244200 396800 244274 396828
rect 40034 396720 40040 396772
rect 40092 396760 40098 396772
rect 212534 396760 212540 396772
rect 40092 396732 212540 396760
rect 40092 396720 40098 396732
rect 212534 396720 212540 396732
rect 212592 396720 212598 396772
rect 212902 396720 212908 396772
rect 212960 396760 212966 396772
rect 213362 396760 213368 396772
rect 212960 396732 213368 396760
rect 212960 396720 212966 396732
rect 213362 396720 213368 396732
rect 213420 396720 213426 396772
rect 214098 396720 214104 396772
rect 214156 396760 214162 396772
rect 214558 396760 214564 396772
rect 214156 396732 214564 396760
rect 214156 396720 214162 396732
rect 214558 396720 214564 396732
rect 214616 396720 214622 396772
rect 226702 396720 226708 396772
rect 226760 396760 226766 396772
rect 227162 396760 227168 396772
rect 226760 396732 227168 396760
rect 226760 396720 226766 396732
rect 227162 396720 227168 396732
rect 227220 396720 227226 396772
rect 229554 396720 229560 396772
rect 229612 396720 229618 396772
rect 231026 396720 231032 396772
rect 231084 396760 231090 396772
rect 231486 396760 231492 396772
rect 231084 396732 231492 396760
rect 231084 396720 231090 396732
rect 231486 396720 231492 396732
rect 231544 396720 231550 396772
rect 232222 396720 232228 396772
rect 232280 396760 232286 396772
rect 232280 396732 232636 396760
rect 232280 396720 232286 396732
rect 209866 396652 209872 396704
rect 209924 396692 209930 396704
rect 210510 396692 210516 396704
rect 209924 396664 210516 396692
rect 209924 396652 209930 396664
rect 210510 396652 210516 396664
rect 210568 396652 210574 396704
rect 211338 396652 211344 396704
rect 211396 396692 211402 396704
rect 212074 396692 212080 396704
rect 211396 396664 212080 396692
rect 211396 396652 211402 396664
rect 212074 396652 212080 396664
rect 212132 396652 212138 396704
rect 212810 396652 212816 396704
rect 212868 396692 212874 396704
rect 213822 396692 213828 396704
rect 212868 396664 213828 396692
rect 212868 396652 212874 396664
rect 213822 396652 213828 396664
rect 213880 396652 213886 396704
rect 214190 396652 214196 396704
rect 214248 396692 214254 396704
rect 214926 396692 214932 396704
rect 214248 396664 214932 396692
rect 214248 396652 214254 396664
rect 214926 396652 214932 396664
rect 214984 396652 214990 396704
rect 225782 396652 225788 396704
rect 225840 396692 225846 396704
rect 226242 396692 226248 396704
rect 225840 396664 226248 396692
rect 225840 396652 225846 396664
rect 226242 396652 226248 396664
rect 226300 396652 226306 396704
rect 227898 396652 227904 396704
rect 227956 396692 227962 396704
rect 228174 396692 228180 396704
rect 227956 396664 228180 396692
rect 227956 396652 227962 396664
rect 228174 396652 228180 396664
rect 228232 396652 228238 396704
rect 228266 396652 228272 396704
rect 228324 396692 228330 396704
rect 228818 396692 228824 396704
rect 228324 396664 228824 396692
rect 228324 396652 228330 396664
rect 228818 396652 228824 396664
rect 228876 396652 228882 396704
rect 209958 396584 209964 396636
rect 210016 396624 210022 396636
rect 210878 396624 210884 396636
rect 210016 396596 210884 396624
rect 210016 396584 210022 396596
rect 210878 396584 210884 396596
rect 210936 396584 210942 396636
rect 211246 396584 211252 396636
rect 211304 396624 211310 396636
rect 211982 396624 211988 396636
rect 211304 396596 211988 396624
rect 211304 396584 211310 396596
rect 211982 396584 211988 396596
rect 212040 396584 212046 396636
rect 212902 396584 212908 396636
rect 212960 396624 212966 396636
rect 213270 396624 213276 396636
rect 212960 396596 213276 396624
rect 212960 396584 212966 396596
rect 213270 396584 213276 396596
rect 213328 396584 213334 396636
rect 214466 396584 214472 396636
rect 214524 396624 214530 396636
rect 214742 396624 214748 396636
rect 214524 396596 214748 396624
rect 214524 396584 214530 396596
rect 214742 396584 214748 396596
rect 214800 396584 214806 396636
rect 211522 396516 211528 396568
rect 211580 396556 211586 396568
rect 212350 396556 212356 396568
rect 211580 396528 212356 396556
rect 211580 396516 211586 396528
rect 212350 396516 212356 396528
rect 212408 396516 212414 396568
rect 212994 396516 213000 396568
rect 213052 396556 213058 396568
rect 213638 396556 213644 396568
rect 213052 396528 213644 396556
rect 213052 396516 213058 396528
rect 213638 396516 213644 396528
rect 213696 396516 213702 396568
rect 214558 396516 214564 396568
rect 214616 396556 214622 396568
rect 215202 396556 215208 396568
rect 214616 396528 215208 396556
rect 214616 396516 214622 396528
rect 215202 396516 215208 396528
rect 215260 396516 215266 396568
rect 226702 396516 226708 396568
rect 226760 396556 226766 396568
rect 227254 396556 227260 396568
rect 226760 396528 227260 396556
rect 226760 396516 226766 396528
rect 227254 396516 227260 396528
rect 227312 396516 227318 396568
rect 227898 396516 227904 396568
rect 227956 396556 227962 396568
rect 228082 396556 228088 396568
rect 227956 396528 228088 396556
rect 227956 396516 227962 396528
rect 228082 396516 228088 396528
rect 228140 396516 228146 396568
rect 229370 396516 229376 396568
rect 229428 396556 229434 396568
rect 229572 396556 229600 396720
rect 232608 396568 232636 396732
rect 232682 396720 232688 396772
rect 232740 396720 232746 396772
rect 234982 396720 234988 396772
rect 235040 396760 235046 396772
rect 235166 396760 235172 396772
rect 235040 396732 235172 396760
rect 235040 396720 235046 396732
rect 235166 396720 235172 396732
rect 235224 396720 235230 396772
rect 235258 396720 235264 396772
rect 235316 396760 235322 396772
rect 235902 396760 235908 396772
rect 235316 396732 235908 396760
rect 235316 396720 235322 396732
rect 235902 396720 235908 396732
rect 235960 396720 235966 396772
rect 236270 396720 236276 396772
rect 236328 396760 236334 396772
rect 237006 396760 237012 396772
rect 236328 396732 237012 396760
rect 236328 396720 236334 396732
rect 237006 396720 237012 396732
rect 237064 396720 237070 396772
rect 237374 396720 237380 396772
rect 237432 396760 237438 396772
rect 237742 396760 237748 396772
rect 237432 396732 237748 396760
rect 237432 396720 237438 396732
rect 237742 396720 237748 396732
rect 237800 396720 237806 396772
rect 238018 396720 238024 396772
rect 238076 396720 238082 396772
rect 240318 396720 240324 396772
rect 240376 396720 240382 396772
rect 240594 396720 240600 396772
rect 240652 396760 240658 396772
rect 240778 396760 240784 396772
rect 240652 396732 240784 396760
rect 240652 396720 240658 396732
rect 240778 396720 240784 396732
rect 240836 396720 240842 396772
rect 241514 396720 241520 396772
rect 241572 396760 241578 396772
rect 241882 396760 241888 396772
rect 241572 396732 241888 396760
rect 241572 396720 241578 396732
rect 241882 396720 241888 396732
rect 241940 396720 241946 396772
rect 243078 396720 243084 396772
rect 243136 396720 243142 396772
rect 243354 396720 243360 396772
rect 243412 396760 243418 396772
rect 243722 396760 243728 396772
rect 243412 396732 243728 396760
rect 243412 396720 243418 396732
rect 243722 396720 243728 396732
rect 243780 396720 243786 396772
rect 244246 396760 244274 396800
rect 249058 396788 249064 396840
rect 249116 396828 249122 396840
rect 402974 396828 402980 396840
rect 249116 396800 402980 396828
rect 249116 396788 249122 396800
rect 402974 396788 402980 396800
rect 403032 396788 403038 396840
rect 409874 396760 409880 396772
rect 244246 396732 409880 396760
rect 409874 396720 409880 396732
rect 409932 396720 409938 396772
rect 229428 396528 229600 396556
rect 229428 396516 229434 396528
rect 232222 396516 232228 396568
rect 232280 396556 232286 396568
rect 232406 396556 232412 396568
rect 232280 396528 232412 396556
rect 232280 396516 232286 396528
rect 232406 396516 232412 396528
rect 232464 396516 232470 396568
rect 232590 396516 232596 396568
rect 232648 396516 232654 396568
rect 212626 396448 212632 396500
rect 212684 396488 212690 396500
rect 213730 396488 213736 396500
rect 212684 396460 213736 396488
rect 212684 396448 212690 396460
rect 213730 396448 213736 396460
rect 213788 396448 213794 396500
rect 226794 396448 226800 396500
rect 226852 396488 226858 396500
rect 227530 396488 227536 396500
rect 226852 396460 227536 396488
rect 226852 396448 226858 396460
rect 227530 396448 227536 396460
rect 227588 396448 227594 396500
rect 229462 396448 229468 396500
rect 229520 396488 229526 396500
rect 229922 396488 229928 396500
rect 229520 396460 229928 396488
rect 229520 396448 229526 396460
rect 229922 396448 229928 396460
rect 229980 396448 229986 396500
rect 210234 396380 210240 396432
rect 210292 396420 210298 396432
rect 210970 396420 210976 396432
rect 210292 396392 210976 396420
rect 210292 396380 210298 396392
rect 210970 396380 210976 396392
rect 211028 396380 211034 396432
rect 228082 396380 228088 396432
rect 228140 396420 228146 396432
rect 228634 396420 228640 396432
rect 228140 396392 228640 396420
rect 228140 396380 228146 396392
rect 228634 396380 228640 396392
rect 228692 396380 228698 396432
rect 229094 396380 229100 396432
rect 229152 396420 229158 396432
rect 229646 396420 229652 396432
rect 229152 396392 229652 396420
rect 229152 396380 229158 396392
rect 229646 396380 229652 396392
rect 229704 396380 229710 396432
rect 230842 396380 230848 396432
rect 230900 396420 230906 396432
rect 231210 396420 231216 396432
rect 230900 396392 231216 396420
rect 230900 396380 230906 396392
rect 231210 396380 231216 396392
rect 231268 396380 231274 396432
rect 232406 396380 232412 396432
rect 232464 396420 232470 396432
rect 232700 396420 232728 396720
rect 236362 396652 236368 396704
rect 236420 396692 236426 396704
rect 236730 396692 236736 396704
rect 236420 396664 236736 396692
rect 236420 396652 236426 396664
rect 236730 396652 236736 396664
rect 236788 396652 236794 396704
rect 233510 396516 233516 396568
rect 233568 396556 233574 396568
rect 233970 396556 233976 396568
rect 233568 396528 233976 396556
rect 233568 396516 233574 396528
rect 233970 396516 233976 396528
rect 234028 396516 234034 396568
rect 234522 396516 234528 396568
rect 234580 396556 234586 396568
rect 235074 396556 235080 396568
rect 234580 396528 235080 396556
rect 234580 396516 234586 396528
rect 235074 396516 235080 396528
rect 235132 396516 235138 396568
rect 237650 396516 237656 396568
rect 237708 396556 237714 396568
rect 238036 396556 238064 396720
rect 239122 396652 239128 396704
rect 239180 396692 239186 396704
rect 239490 396692 239496 396704
rect 239180 396664 239496 396692
rect 239180 396652 239186 396664
rect 239490 396652 239496 396664
rect 239548 396652 239554 396704
rect 237708 396528 238064 396556
rect 237708 396516 237714 396528
rect 239030 396516 239036 396568
rect 239088 396556 239094 396568
rect 239582 396556 239588 396568
rect 239088 396528 239588 396556
rect 239088 396516 239094 396528
rect 239582 396516 239588 396528
rect 239640 396516 239646 396568
rect 240336 396556 240364 396720
rect 240686 396556 240692 396568
rect 240336 396528 240692 396556
rect 240686 396516 240692 396528
rect 240744 396516 240750 396568
rect 243096 396556 243124 396720
rect 243446 396556 243452 396568
rect 243096 396528 243452 396556
rect 243446 396516 243452 396528
rect 243504 396516 243510 396568
rect 234798 396448 234804 396500
rect 234856 396488 234862 396500
rect 235534 396488 235540 396500
rect 234856 396460 235540 396488
rect 234856 396448 234862 396460
rect 235534 396448 235540 396460
rect 235592 396448 235598 396500
rect 237926 396448 237932 396500
rect 237984 396488 237990 396500
rect 238110 396488 238116 396500
rect 237984 396460 238116 396488
rect 237984 396448 237990 396460
rect 238110 396448 238116 396460
rect 238168 396448 238174 396500
rect 240134 396448 240140 396500
rect 240192 396488 240198 396500
rect 240410 396488 240416 396500
rect 240192 396460 240416 396488
rect 240192 396448 240198 396460
rect 240410 396448 240416 396460
rect 240468 396448 240474 396500
rect 240502 396448 240508 396500
rect 240560 396488 240566 396500
rect 241146 396488 241152 396500
rect 240560 396460 241152 396488
rect 240560 396448 240566 396460
rect 241146 396448 241152 396460
rect 241204 396448 241210 396500
rect 242894 396448 242900 396500
rect 242952 396488 242958 396500
rect 243262 396488 243268 396500
rect 242952 396460 243268 396488
rect 242952 396448 242958 396460
rect 243262 396448 243268 396460
rect 243320 396448 243326 396500
rect 232464 396392 232728 396420
rect 232464 396380 232470 396392
rect 233326 396380 233332 396432
rect 233384 396420 233390 396432
rect 233878 396420 233884 396432
rect 233384 396392 233884 396420
rect 233384 396380 233390 396392
rect 233878 396380 233884 396392
rect 233936 396380 233942 396432
rect 236086 396380 236092 396432
rect 236144 396420 236150 396432
rect 236638 396420 236644 396432
rect 236144 396392 236644 396420
rect 236144 396380 236150 396392
rect 236638 396380 236644 396392
rect 236696 396380 236702 396432
rect 237834 396380 237840 396432
rect 237892 396420 237898 396432
rect 238202 396420 238208 396432
rect 237892 396392 238208 396420
rect 237892 396380 237898 396392
rect 238202 396380 238208 396392
rect 238260 396380 238266 396432
rect 240318 396380 240324 396432
rect 240376 396420 240382 396432
rect 241054 396420 241060 396432
rect 240376 396392 241060 396420
rect 240376 396380 240382 396392
rect 241054 396380 241060 396392
rect 241112 396380 241118 396432
rect 241698 396380 241704 396432
rect 241756 396420 241762 396432
rect 241974 396420 241980 396432
rect 241756 396392 241980 396420
rect 241756 396380 241762 396392
rect 241974 396380 241980 396392
rect 242032 396380 242038 396432
rect 243170 396380 243176 396432
rect 243228 396420 243234 396432
rect 243814 396420 243820 396432
rect 243228 396392 243820 396420
rect 243228 396380 243234 396392
rect 243814 396380 243820 396392
rect 243872 396380 243878 396432
rect 210326 396312 210332 396364
rect 210384 396352 210390 396364
rect 211062 396352 211068 396364
rect 210384 396324 211068 396352
rect 210384 396312 210390 396324
rect 211062 396312 211068 396324
rect 211120 396312 211126 396364
rect 222746 396312 222752 396364
rect 222804 396352 222810 396364
rect 227346 396352 227352 396364
rect 222804 396324 227352 396352
rect 222804 396312 222810 396324
rect 227346 396312 227352 396324
rect 227404 396312 227410 396364
rect 230934 396312 230940 396364
rect 230992 396352 230998 396364
rect 231394 396352 231400 396364
rect 230992 396324 231400 396352
rect 230992 396312 230998 396324
rect 231394 396312 231400 396324
rect 231452 396312 231458 396364
rect 233234 396312 233240 396364
rect 233292 396352 233298 396364
rect 233970 396352 233976 396364
rect 233292 396324 233976 396352
rect 233292 396312 233298 396324
rect 233970 396312 233976 396324
rect 234028 396312 234034 396364
rect 235994 396312 236000 396364
rect 236052 396352 236058 396364
rect 236914 396352 236920 396364
rect 236052 396324 236920 396352
rect 236052 396312 236058 396324
rect 236914 396312 236920 396324
rect 236972 396312 236978 396364
rect 237558 396312 237564 396364
rect 237616 396352 237622 396364
rect 237926 396352 237932 396364
rect 237616 396324 237932 396352
rect 237616 396312 237622 396324
rect 237926 396312 237932 396324
rect 237984 396312 237990 396364
rect 240410 396312 240416 396364
rect 240468 396352 240474 396364
rect 241238 396352 241244 396364
rect 240468 396324 241244 396352
rect 240468 396312 240474 396324
rect 241238 396312 241244 396324
rect 241296 396312 241302 396364
rect 241606 396312 241612 396364
rect 241664 396352 241670 396364
rect 242158 396352 242164 396364
rect 241664 396324 242164 396352
rect 241664 396312 241670 396324
rect 242158 396312 242164 396324
rect 242216 396312 242222 396364
rect 233878 396244 233884 396296
rect 233936 396284 233942 396296
rect 234062 396284 234068 396296
rect 233936 396256 234068 396284
rect 233936 396244 233942 396256
rect 234062 396244 234068 396256
rect 234120 396244 234126 396296
rect 233234 396176 233240 396228
rect 233292 396216 233298 396228
rect 234154 396216 234160 396228
rect 233292 396188 234160 396216
rect 233292 396176 233298 396188
rect 234154 396176 234160 396188
rect 234212 396176 234218 396228
rect 210510 396108 210516 396160
rect 210568 396148 210574 396160
rect 217226 396148 217232 396160
rect 210568 396120 217232 396148
rect 210568 396108 210574 396120
rect 217226 396108 217232 396120
rect 217284 396108 217290 396160
rect 237650 396108 237656 396160
rect 237708 396148 237714 396160
rect 238294 396148 238300 396160
rect 237708 396120 238300 396148
rect 237708 396108 237714 396120
rect 238294 396108 238300 396120
rect 238352 396108 238358 396160
rect 244182 396108 244188 396160
rect 244240 396148 244246 396160
rect 245470 396148 245476 396160
rect 244240 396120 245476 396148
rect 244240 396108 244246 396120
rect 245470 396108 245476 396120
rect 245528 396108 245534 396160
rect 250438 395972 250444 396024
rect 250496 396012 250502 396024
rect 250806 396012 250812 396024
rect 250496 395984 250812 396012
rect 250496 395972 250502 395984
rect 250806 395972 250812 395984
rect 250864 395972 250870 396024
rect 213178 395904 213184 395956
rect 213236 395944 213242 395956
rect 213454 395944 213460 395956
rect 213236 395916 213460 395944
rect 213236 395904 213242 395916
rect 213454 395904 213460 395916
rect 213512 395904 213518 395956
rect 214006 395904 214012 395956
rect 214064 395944 214070 395956
rect 214374 395944 214380 395956
rect 214064 395916 214380 395944
rect 214064 395904 214070 395916
rect 214374 395904 214380 395916
rect 214432 395904 214438 395956
rect 231578 395904 231584 395956
rect 231636 395944 231642 395956
rect 256234 395944 256240 395956
rect 231636 395916 256240 395944
rect 231636 395904 231642 395916
rect 256234 395904 256240 395916
rect 256292 395904 256298 395956
rect 231486 395836 231492 395888
rect 231544 395876 231550 395888
rect 266354 395876 266360 395888
rect 231544 395848 266360 395876
rect 231544 395836 231550 395848
rect 266354 395836 266360 395848
rect 266412 395836 266418 395888
rect 214006 395768 214012 395820
rect 214064 395808 214070 395820
rect 214834 395808 214840 395820
rect 214064 395780 214840 395808
rect 214064 395768 214070 395780
rect 214834 395768 214840 395780
rect 214892 395768 214898 395820
rect 231302 395768 231308 395820
rect 231360 395808 231366 395820
rect 269114 395808 269120 395820
rect 231360 395780 269120 395808
rect 231360 395768 231366 395780
rect 269114 395768 269120 395780
rect 269172 395768 269178 395820
rect 232866 395700 232872 395752
rect 232924 395740 232930 395752
rect 276014 395740 276020 395752
rect 232924 395712 276020 395740
rect 232924 395700 232930 395712
rect 276014 395700 276020 395712
rect 276072 395700 276078 395752
rect 141418 395632 141424 395684
rect 141476 395672 141482 395684
rect 217502 395672 217508 395684
rect 141476 395644 217508 395672
rect 141476 395632 141482 395644
rect 217502 395632 217508 395644
rect 217560 395632 217566 395684
rect 240042 395632 240048 395684
rect 240100 395672 240106 395684
rect 333974 395672 333980 395684
rect 240100 395644 333980 395672
rect 240100 395632 240106 395644
rect 333974 395632 333980 395644
rect 334032 395632 334038 395684
rect 115934 395564 115940 395616
rect 115992 395604 115998 395616
rect 219342 395604 219348 395616
rect 115992 395576 219348 395604
rect 115992 395564 115998 395576
rect 219342 395564 219348 395576
rect 219400 395564 219406 395616
rect 247310 395564 247316 395616
rect 247368 395604 247374 395616
rect 247678 395604 247684 395616
rect 247368 395576 247684 395604
rect 247368 395564 247374 395576
rect 247678 395564 247684 395576
rect 247736 395564 247742 395616
rect 250162 395564 250168 395616
rect 250220 395604 250226 395616
rect 250438 395604 250444 395616
rect 250220 395576 250444 395604
rect 250220 395564 250226 395576
rect 250438 395564 250444 395576
rect 250496 395564 250502 395616
rect 252002 395564 252008 395616
rect 252060 395604 252066 395616
rect 535454 395604 535460 395616
rect 252060 395576 535460 395604
rect 252060 395564 252066 395576
rect 535454 395564 535460 395576
rect 535512 395564 535518 395616
rect 77294 395496 77300 395548
rect 77352 395536 77358 395548
rect 216398 395536 216404 395548
rect 77352 395508 216404 395536
rect 77352 395496 77358 395508
rect 216398 395496 216404 395508
rect 216456 395496 216462 395548
rect 253106 395496 253112 395548
rect 253164 395536 253170 395548
rect 549254 395536 549260 395548
rect 253164 395508 549260 395536
rect 253164 395496 253170 395508
rect 549254 395496 549260 395508
rect 549312 395496 549318 395548
rect 52454 395428 52460 395480
rect 52512 395468 52518 395480
rect 214374 395468 214380 395480
rect 52512 395440 214380 395468
rect 52512 395428 52518 395440
rect 214374 395428 214380 395440
rect 214432 395428 214438 395480
rect 253934 395428 253940 395480
rect 253992 395468 253998 395480
rect 560294 395468 560300 395480
rect 253992 395440 560300 395468
rect 253992 395428 253998 395440
rect 560294 395428 560300 395440
rect 560352 395428 560358 395480
rect 30374 395360 30380 395412
rect 30432 395400 30438 395412
rect 212534 395400 212540 395412
rect 30432 395372 212540 395400
rect 30432 395360 30438 395372
rect 212534 395360 212540 395372
rect 212592 395360 212598 395412
rect 254210 395360 254216 395412
rect 254268 395400 254274 395412
rect 564526 395400 564532 395412
rect 254268 395372 564532 395400
rect 254268 395360 254274 395372
rect 564526 395360 564532 395372
rect 564584 395360 564590 395412
rect 27614 395292 27620 395344
rect 27672 395332 27678 395344
rect 212166 395332 212172 395344
rect 27672 395304 212172 395332
rect 27672 395292 27678 395304
rect 212166 395292 212172 395304
rect 212224 395292 212230 395344
rect 226518 395292 226524 395344
rect 226576 395332 226582 395344
rect 226886 395332 226892 395344
rect 226576 395304 226892 395332
rect 226576 395292 226582 395304
rect 226886 395292 226892 395304
rect 226944 395292 226950 395344
rect 254762 395292 254768 395344
rect 254820 395332 254826 395344
rect 571334 395332 571340 395344
rect 254820 395304 571340 395332
rect 254820 395292 254826 395304
rect 571334 395292 571340 395304
rect 571392 395292 571398 395344
rect 214374 395156 214380 395208
rect 214432 395196 214438 395208
rect 214650 395196 214656 395208
rect 214432 395168 214656 395196
rect 214432 395156 214438 395168
rect 214650 395156 214656 395168
rect 214708 395156 214714 395208
rect 251542 395020 251548 395072
rect 251600 395060 251606 395072
rect 252002 395060 252008 395072
rect 251600 395032 252008 395060
rect 251600 395020 251606 395032
rect 252002 395020 252008 395032
rect 252060 395020 252066 395072
rect 216398 394680 216404 394732
rect 216456 394720 216462 394732
rect 223298 394720 223304 394732
rect 216456 394692 223304 394720
rect 216456 394680 216462 394692
rect 223298 394680 223304 394692
rect 223356 394680 223362 394732
rect 228358 394680 228364 394732
rect 228416 394720 228422 394732
rect 231118 394720 231124 394732
rect 228416 394692 231124 394720
rect 228416 394680 228422 394692
rect 231118 394680 231124 394692
rect 231176 394680 231182 394732
rect 254026 394680 254032 394732
rect 254084 394720 254090 394732
rect 254394 394720 254400 394732
rect 254084 394692 254400 394720
rect 254084 394680 254090 394692
rect 254394 394680 254400 394692
rect 254452 394680 254458 394732
rect 215294 394612 215300 394664
rect 215352 394652 215358 394664
rect 218882 394652 218888 394664
rect 215352 394624 218888 394652
rect 215352 394612 215358 394624
rect 218882 394612 218888 394624
rect 218940 394612 218946 394664
rect 225598 394612 225604 394664
rect 225656 394652 225662 394664
rect 227070 394652 227076 394664
rect 225656 394624 227076 394652
rect 225656 394612 225662 394624
rect 227070 394612 227076 394624
rect 227128 394612 227134 394664
rect 244550 394612 244556 394664
rect 244608 394652 244614 394664
rect 245562 394652 245568 394664
rect 244608 394624 245568 394652
rect 244608 394612 244614 394624
rect 245562 394612 245568 394624
rect 245620 394612 245626 394664
rect 247954 394612 247960 394664
rect 248012 394652 248018 394664
rect 258718 394652 258724 394664
rect 248012 394624 258724 394652
rect 248012 394612 248018 394624
rect 258718 394612 258724 394624
rect 258776 394612 258782 394664
rect 215386 394544 215392 394596
rect 215444 394584 215450 394596
rect 215938 394584 215944 394596
rect 215444 394556 215944 394584
rect 215444 394544 215450 394556
rect 215938 394544 215944 394556
rect 215996 394544 216002 394596
rect 251266 394544 251272 394596
rect 251324 394584 251330 394596
rect 251818 394584 251824 394596
rect 251324 394556 251824 394584
rect 251324 394544 251330 394556
rect 251818 394544 251824 394556
rect 251876 394544 251882 394596
rect 253934 394544 253940 394596
rect 253992 394584 253998 394596
rect 254578 394584 254584 394596
rect 253992 394556 254584 394584
rect 253992 394544 253998 394556
rect 254578 394544 254584 394556
rect 254636 394544 254642 394596
rect 224494 394516 224500 394528
rect 215266 394488 224500 394516
rect 4154 394408 4160 394460
rect 4212 394448 4218 394460
rect 209774 394448 209780 394460
rect 4212 394420 209780 394448
rect 4212 394408 4218 394420
rect 209774 394408 209780 394420
rect 209832 394408 209838 394460
rect 209130 394340 209136 394392
rect 209188 394380 209194 394392
rect 215266 394380 215294 394488
rect 224494 394476 224500 394488
rect 224552 394476 224558 394528
rect 234338 394476 234344 394528
rect 234396 394516 234402 394528
rect 304994 394516 305000 394528
rect 234396 394488 305000 394516
rect 234396 394476 234402 394488
rect 304994 394476 305000 394488
rect 305052 394476 305058 394528
rect 235626 394408 235632 394460
rect 235684 394448 235690 394460
rect 322934 394448 322940 394460
rect 235684 394420 322940 394448
rect 235684 394408 235690 394420
rect 322934 394408 322940 394420
rect 322992 394408 322998 394460
rect 224218 394380 224224 394392
rect 209188 394352 215294 394380
rect 215404 394352 224224 394380
rect 209188 394340 209194 394352
rect 189074 394272 189080 394324
rect 189132 394312 189138 394324
rect 212442 394312 212448 394324
rect 189132 394284 212448 394312
rect 189132 394272 189138 394284
rect 212442 394272 212448 394284
rect 212500 394272 212506 394324
rect 178034 394204 178040 394256
rect 178092 394244 178098 394256
rect 215404 394244 215432 394352
rect 224218 394340 224224 394352
rect 224276 394340 224282 394392
rect 237006 394340 237012 394392
rect 237064 394380 237070 394392
rect 332594 394380 332600 394392
rect 237064 394352 332600 394380
rect 237064 394340 237070 394352
rect 332594 394340 332600 394352
rect 332652 394340 332658 394392
rect 221090 394272 221096 394324
rect 221148 394312 221154 394324
rect 221550 394312 221556 394324
rect 221148 394284 221556 394312
rect 221148 394272 221154 394284
rect 221550 394272 221556 394284
rect 221608 394272 221614 394324
rect 223758 394272 223764 394324
rect 223816 394312 223822 394324
rect 224310 394312 224316 394324
rect 223816 394284 224316 394312
rect 223816 394272 223822 394284
rect 224310 394272 224316 394284
rect 224368 394272 224374 394324
rect 236822 394272 236828 394324
rect 236880 394312 236886 394324
rect 340874 394312 340880 394324
rect 236880 394284 340880 394312
rect 236880 394272 236886 394284
rect 340874 394272 340880 394284
rect 340932 394272 340938 394324
rect 220446 394244 220452 394256
rect 178092 394216 215432 394244
rect 215496 394216 220452 394244
rect 178092 394204 178098 394216
rect 133874 394136 133880 394188
rect 133932 394176 133938 394188
rect 215294 394176 215300 394188
rect 133932 394148 215300 394176
rect 133932 394136 133938 394148
rect 215294 394136 215300 394148
rect 215352 394136 215358 394188
rect 129734 394068 129740 394120
rect 129792 394108 129798 394120
rect 215496 394108 215524 394216
rect 220446 394204 220452 394216
rect 220504 394204 220510 394256
rect 238386 394204 238392 394256
rect 238444 394244 238450 394256
rect 347774 394244 347780 394256
rect 238444 394216 347780 394244
rect 238444 394204 238450 394216
rect 347774 394204 347780 394216
rect 347832 394204 347838 394256
rect 215570 394136 215576 394188
rect 215628 394176 215634 394188
rect 216214 394176 216220 394188
rect 215628 394148 216220 394176
rect 215628 394136 215634 394148
rect 216214 394136 216220 394148
rect 216272 394136 216278 394188
rect 216950 394136 216956 394188
rect 217008 394176 217014 394188
rect 217410 394176 217416 394188
rect 217008 394148 217416 394176
rect 217008 394136 217014 394148
rect 217410 394136 217416 394148
rect 217468 394136 217474 394188
rect 220906 394136 220912 394188
rect 220964 394176 220970 394188
rect 222010 394176 222016 394188
rect 220964 394148 222016 394176
rect 220964 394136 220970 394148
rect 222010 394136 222016 394148
rect 222068 394136 222074 394188
rect 222378 394136 222384 394188
rect 222436 394176 222442 394188
rect 222930 394176 222936 394188
rect 222436 394148 222936 394176
rect 222436 394136 222442 394148
rect 222930 394136 222936 394148
rect 222988 394136 222994 394188
rect 223850 394136 223856 394188
rect 223908 394176 223914 394188
rect 224586 394176 224592 394188
rect 223908 394148 224592 394176
rect 223908 394136 223914 394148
rect 224586 394136 224592 394148
rect 224644 394136 224650 394188
rect 243998 394136 244004 394188
rect 244056 394176 244062 394188
rect 365714 394176 365720 394188
rect 244056 394148 365720 394176
rect 244056 394136 244062 394148
rect 365714 394136 365720 394148
rect 365772 394136 365778 394188
rect 217686 394108 217692 394120
rect 129792 394080 215524 394108
rect 215588 394080 217692 394108
rect 129792 394068 129798 394080
rect 92474 394000 92480 394052
rect 92532 394040 92538 394052
rect 215588 394040 215616 394080
rect 217686 394068 217692 394080
rect 217744 394068 217750 394120
rect 218238 394068 218244 394120
rect 218296 394108 218302 394120
rect 218974 394108 218980 394120
rect 218296 394080 218980 394108
rect 218296 394068 218302 394080
rect 218974 394068 218980 394080
rect 219032 394068 219038 394120
rect 219526 394068 219532 394120
rect 219584 394108 219590 394120
rect 220354 394108 220360 394120
rect 219584 394080 220360 394108
rect 219584 394068 219590 394080
rect 220354 394068 220360 394080
rect 220412 394068 220418 394120
rect 221182 394068 221188 394120
rect 221240 394108 221246 394120
rect 221826 394108 221832 394120
rect 221240 394080 221832 394108
rect 221240 394068 221246 394080
rect 221826 394068 221832 394080
rect 221884 394068 221890 394120
rect 223942 394068 223948 394120
rect 224000 394108 224006 394120
rect 224862 394108 224868 394120
rect 224000 394080 224868 394108
rect 224000 394068 224006 394080
rect 224862 394068 224868 394080
rect 224920 394068 224926 394120
rect 240226 394068 240232 394120
rect 240284 394108 240290 394120
rect 382274 394108 382280 394120
rect 240284 394080 382280 394108
rect 240284 394068 240290 394080
rect 382274 394068 382280 394080
rect 382332 394068 382338 394120
rect 92532 394012 215616 394040
rect 92532 394000 92538 394012
rect 215662 394000 215668 394052
rect 215720 394040 215726 394052
rect 216214 394040 216220 394052
rect 215720 394012 216220 394040
rect 215720 394000 215726 394012
rect 216214 394000 216220 394012
rect 216272 394000 216278 394052
rect 216858 394000 216864 394052
rect 216916 394040 216922 394052
rect 217870 394040 217876 394052
rect 216916 394012 217876 394040
rect 216916 394000 216922 394012
rect 217870 394000 217876 394012
rect 217928 394000 217934 394052
rect 218606 394000 218612 394052
rect 218664 394040 218670 394052
rect 219066 394040 219072 394052
rect 218664 394012 219072 394040
rect 218664 394000 218670 394012
rect 219066 394000 219072 394012
rect 219124 394000 219130 394052
rect 219802 394000 219808 394052
rect 219860 394040 219866 394052
rect 220262 394040 220268 394052
rect 219860 394012 220268 394040
rect 219860 394000 219866 394012
rect 220262 394000 220268 394012
rect 220320 394000 220326 394052
rect 221550 394000 221556 394052
rect 221608 394040 221614 394052
rect 221918 394040 221924 394052
rect 221608 394012 221924 394040
rect 221608 394000 221614 394012
rect 221918 394000 221924 394012
rect 221976 394000 221982 394052
rect 224310 394000 224316 394052
rect 224368 394040 224374 394052
rect 224770 394040 224776 394052
rect 224368 394012 224776 394040
rect 224368 394000 224374 394012
rect 224770 394000 224776 394012
rect 224828 394000 224834 394052
rect 225046 394040 225052 394052
rect 224926 394012 225052 394040
rect 210418 393932 210424 393984
rect 210476 393972 210482 393984
rect 224926 393972 224954 394012
rect 225046 394000 225052 394012
rect 225104 394000 225110 394052
rect 244918 394000 244924 394052
rect 244976 394000 244982 394052
rect 252738 394000 252744 394052
rect 252796 394040 252802 394052
rect 253106 394040 253112 394052
rect 252796 394012 253112 394040
rect 252796 394000 252802 394012
rect 253106 394000 253112 394012
rect 253164 394000 253170 394052
rect 440234 394040 440240 394052
rect 253308 394012 440240 394040
rect 210476 393944 224954 393972
rect 210476 393932 210482 393944
rect 209774 393864 209780 393916
rect 209832 393904 209838 393916
rect 210510 393904 210516 393916
rect 209832 393876 210516 393904
rect 209832 393864 209838 393876
rect 210510 393864 210516 393876
rect 210568 393864 210574 393916
rect 215662 393864 215668 393916
rect 215720 393904 215726 393916
rect 216306 393904 216312 393916
rect 215720 393876 216312 393904
rect 215720 393864 215726 393876
rect 216306 393864 216312 393876
rect 216364 393864 216370 393916
rect 218422 393864 218428 393916
rect 218480 393904 218486 393916
rect 218790 393904 218796 393916
rect 218480 393876 218796 393904
rect 218480 393864 218486 393876
rect 218790 393864 218796 393876
rect 218848 393864 218854 393916
rect 219710 393864 219716 393916
rect 219768 393904 219774 393916
rect 220170 393904 220176 393916
rect 219768 393876 220176 393904
rect 219768 393864 219774 393876
rect 220170 393864 220176 393876
rect 220228 393864 220234 393916
rect 221366 393864 221372 393916
rect 221424 393904 221430 393916
rect 221734 393904 221740 393916
rect 221424 393876 221740 393904
rect 221424 393864 221430 393876
rect 221734 393864 221740 393876
rect 221792 393864 221798 393916
rect 222470 393864 222476 393916
rect 222528 393904 222534 393916
rect 222930 393904 222936 393916
rect 222528 393876 222936 393904
rect 222528 393864 222534 393876
rect 222930 393864 222936 393876
rect 222988 393864 222994 393916
rect 224034 393864 224040 393916
rect 224092 393904 224098 393916
rect 224402 393904 224408 393916
rect 224092 393876 224408 393904
rect 224092 393864 224098 393876
rect 224402 393864 224408 393876
rect 224460 393864 224466 393916
rect 216030 393796 216036 393848
rect 216088 393836 216094 393848
rect 216582 393836 216588 393848
rect 216088 393808 216588 393836
rect 216088 393796 216094 393808
rect 216582 393796 216588 393808
rect 216640 393796 216646 393848
rect 218330 393796 218336 393848
rect 218388 393836 218394 393848
rect 219250 393836 219256 393848
rect 218388 393808 219256 393836
rect 218388 393796 218394 393808
rect 219250 393796 219256 393808
rect 219308 393796 219314 393848
rect 219618 393796 219624 393848
rect 219676 393836 219682 393848
rect 220630 393836 220636 393848
rect 219676 393808 220636 393836
rect 219676 393796 219682 393808
rect 220630 393796 220636 393808
rect 220688 393796 220694 393848
rect 220998 393796 221004 393848
rect 221056 393836 221062 393848
rect 222102 393836 222108 393848
rect 221056 393808 222108 393836
rect 221056 393796 221062 393808
rect 222102 393796 222108 393808
rect 222160 393796 222166 393848
rect 244458 393796 244464 393848
rect 244516 393836 244522 393848
rect 244936 393836 244964 394000
rect 246298 393932 246304 393984
rect 246356 393972 246362 393984
rect 246942 393972 246948 393984
rect 246356 393944 246948 393972
rect 246356 393932 246362 393944
rect 246942 393932 246948 393944
rect 247000 393932 247006 393984
rect 251358 393932 251364 393984
rect 251416 393972 251422 393984
rect 251542 393972 251548 393984
rect 251416 393944 251548 393972
rect 251416 393932 251422 393944
rect 251542 393932 251548 393944
rect 251600 393932 251606 393984
rect 245562 393864 245568 393916
rect 245620 393904 245626 393916
rect 253308 393904 253336 394012
rect 440234 394000 440240 394012
rect 440292 394000 440298 394052
rect 492674 393972 492680 393984
rect 245620 393876 253336 393904
rect 253906 393944 492680 393972
rect 245620 393864 245626 393876
rect 244516 393808 244964 393836
rect 244516 393796 244522 393808
rect 245838 393796 245844 393848
rect 245896 393836 245902 393848
rect 246574 393836 246580 393848
rect 245896 393808 246580 393836
rect 245896 393796 245902 393808
rect 246574 393796 246580 393808
rect 246632 393796 246638 393848
rect 250070 393796 250076 393848
rect 250128 393836 250134 393848
rect 250254 393836 250260 393848
rect 250128 393808 250260 393836
rect 250128 393796 250134 393808
rect 250254 393796 250260 393808
rect 250312 393796 250318 393848
rect 251174 393796 251180 393848
rect 251232 393836 251238 393848
rect 251358 393836 251364 393848
rect 251232 393808 251364 393836
rect 251232 393796 251238 393808
rect 251358 393796 251364 393808
rect 251416 393796 251422 393848
rect 251634 393796 251640 393848
rect 251692 393836 251698 393848
rect 251910 393836 251916 393848
rect 251692 393808 251916 393836
rect 251692 393796 251698 393808
rect 251910 393796 251916 393808
rect 251968 393796 251974 393848
rect 252830 393796 252836 393848
rect 252888 393836 252894 393848
rect 253198 393836 253204 393848
rect 252888 393808 253204 393836
rect 252888 393796 252894 393808
rect 253198 393796 253204 393808
rect 253256 393796 253262 393848
rect 215478 393728 215484 393780
rect 215536 393768 215542 393780
rect 216490 393768 216496 393780
rect 215536 393740 216496 393768
rect 215536 393728 215542 393740
rect 216490 393728 216496 393740
rect 216548 393728 216554 393780
rect 218422 393728 218428 393780
rect 218480 393768 218486 393780
rect 219158 393768 219164 393780
rect 218480 393740 219164 393768
rect 218480 393728 218486 393740
rect 219158 393728 219164 393740
rect 219216 393728 219222 393780
rect 244366 393728 244372 393780
rect 244424 393768 244430 393780
rect 245194 393768 245200 393780
rect 244424 393740 245200 393768
rect 244424 393728 244430 393740
rect 245194 393728 245200 393740
rect 245252 393728 245258 393780
rect 247218 393728 247224 393780
rect 247276 393768 247282 393780
rect 247276 393740 247356 393768
rect 247276 393728 247282 393740
rect 215938 393660 215944 393712
rect 215996 393700 216002 393712
rect 216398 393700 216404 393712
rect 215996 393672 216404 393700
rect 215996 393660 216002 393672
rect 216398 393660 216404 393672
rect 216456 393660 216462 393712
rect 247328 393576 247356 393740
rect 252738 393728 252744 393780
rect 252796 393768 252802 393780
rect 253474 393768 253480 393780
rect 252796 393740 253480 393768
rect 252796 393728 252802 393740
rect 253474 393728 253480 393740
rect 253532 393728 253538 393780
rect 251174 393660 251180 393712
rect 251232 393700 251238 393712
rect 252094 393700 252100 393712
rect 251232 393672 252100 393700
rect 251232 393660 251238 393672
rect 252094 393660 252100 393672
rect 252152 393660 252158 393712
rect 252646 393660 252652 393712
rect 252704 393700 252710 393712
rect 252922 393700 252928 393712
rect 252704 393672 252928 393700
rect 252704 393660 252710 393672
rect 252922 393660 252928 393672
rect 252980 393660 252986 393712
rect 248690 393592 248696 393644
rect 248748 393632 248754 393644
rect 253906 393632 253934 393944
rect 492674 393932 492680 393944
rect 492732 393932 492738 393984
rect 254118 393864 254124 393916
rect 254176 393904 254182 393916
rect 254854 393904 254860 393916
rect 254176 393876 254860 393904
rect 254176 393864 254182 393876
rect 254854 393864 254860 393876
rect 254912 393864 254918 393916
rect 248748 393604 253934 393632
rect 248748 393592 248754 393604
rect 247310 393524 247316 393576
rect 247368 393524 247374 393576
rect 252922 393252 252928 393304
rect 252980 393292 252986 393304
rect 253382 393292 253388 393304
rect 252980 393264 253388 393292
rect 252980 393252 252986 393264
rect 253382 393252 253388 393264
rect 253440 393252 253446 393304
rect 244734 393116 244740 393168
rect 244792 393156 244798 393168
rect 245102 393156 245108 393168
rect 244792 393128 245108 393156
rect 244792 393116 244798 393128
rect 245102 393116 245108 393128
rect 245160 393116 245166 393168
rect 244642 393048 244648 393100
rect 244700 393088 244706 393100
rect 245286 393088 245292 393100
rect 244700 393060 245292 393088
rect 244700 393048 244706 393060
rect 245286 393048 245292 393060
rect 245344 393048 245350 393100
rect 247678 393048 247684 393100
rect 247736 393088 247742 393100
rect 253658 393088 253664 393100
rect 247736 393060 253664 393088
rect 247736 393048 247742 393060
rect 253658 393048 253664 393060
rect 253716 393048 253722 393100
rect 252554 392980 252560 393032
rect 252612 393020 252618 393032
rect 253198 393020 253204 393032
rect 252612 392992 253204 393020
rect 252612 392980 252618 392992
rect 253198 392980 253204 392992
rect 253256 392980 253262 393032
rect 231026 392912 231032 392964
rect 231084 392952 231090 392964
rect 267734 392952 267740 392964
rect 231084 392924 267740 392952
rect 231084 392912 231090 392924
rect 267734 392912 267740 392924
rect 267792 392912 267798 392964
rect 239582 392844 239588 392896
rect 239640 392884 239646 392896
rect 295334 392884 295340 392896
rect 239640 392856 295340 392884
rect 239640 392844 239646 392856
rect 295334 392844 295340 392856
rect 295392 392844 295398 392896
rect 241790 392776 241796 392828
rect 241848 392816 241854 392828
rect 401594 392816 401600 392828
rect 241848 392788 401600 392816
rect 241848 392776 241854 392788
rect 401594 392776 401600 392788
rect 401652 392776 401658 392828
rect 202874 392708 202880 392760
rect 202932 392748 202938 392760
rect 225874 392748 225880 392760
rect 202932 392720 225880 392748
rect 202932 392708 202938 392720
rect 225874 392708 225880 392720
rect 225932 392708 225938 392760
rect 252554 392708 252560 392760
rect 252612 392748 252618 392760
rect 253566 392748 253572 392760
rect 252612 392720 253572 392748
rect 252612 392708 252618 392720
rect 253566 392708 253572 392720
rect 253624 392708 253630 392760
rect 253658 392708 253664 392760
rect 253716 392748 253722 392760
rect 483014 392748 483020 392760
rect 253716 392720 483020 392748
rect 253716 392708 253722 392720
rect 483014 392708 483020 392720
rect 483072 392708 483078 392760
rect 160186 392640 160192 392692
rect 160244 392680 160250 392692
rect 217042 392680 217048 392692
rect 160244 392652 217048 392680
rect 160244 392640 160250 392652
rect 217042 392640 217048 392652
rect 217100 392640 217106 392692
rect 248506 392640 248512 392692
rect 248564 392680 248570 392692
rect 498194 392680 498200 392692
rect 248564 392652 498200 392680
rect 248564 392640 248570 392652
rect 498194 392640 498200 392652
rect 498252 392640 498258 392692
rect 109034 392572 109040 392624
rect 109092 392612 109098 392624
rect 214650 392612 214656 392624
rect 109092 392584 214656 392612
rect 109092 392572 109098 392584
rect 214650 392572 214656 392584
rect 214708 392572 214714 392624
rect 250438 392572 250444 392624
rect 250496 392612 250502 392624
rect 511994 392612 512000 392624
rect 250496 392584 512000 392612
rect 250496 392572 250502 392584
rect 511994 392572 512000 392584
rect 512052 392572 512058 392624
rect 245654 392368 245660 392420
rect 245712 392408 245718 392420
rect 246022 392408 246028 392420
rect 245712 392380 246028 392408
rect 245712 392368 245718 392380
rect 246022 392368 246028 392380
rect 246080 392368 246086 392420
rect 217134 392164 217140 392216
rect 217192 392204 217198 392216
rect 217962 392204 217968 392216
rect 217192 392176 217968 392204
rect 217192 392164 217198 392176
rect 217962 392164 217968 392176
rect 218020 392164 218026 392216
rect 248782 392164 248788 392216
rect 248840 392204 248846 392216
rect 249426 392204 249432 392216
rect 248840 392176 249432 392204
rect 248840 392164 248846 392176
rect 249426 392164 249432 392176
rect 249484 392164 249490 392216
rect 249978 392164 249984 392216
rect 250036 392204 250042 392216
rect 250530 392204 250536 392216
rect 250036 392176 250536 392204
rect 250036 392164 250042 392176
rect 250530 392164 250536 392176
rect 250588 392164 250594 392216
rect 247770 392136 247776 392148
rect 247144 392108 247776 392136
rect 247144 392080 247172 392108
rect 247770 392096 247776 392108
rect 247828 392096 247834 392148
rect 224218 392028 224224 392080
rect 224276 392068 224282 392080
rect 224678 392068 224684 392080
rect 224276 392040 224684 392068
rect 224276 392028 224282 392040
rect 224678 392028 224684 392040
rect 224736 392028 224742 392080
rect 247126 392028 247132 392080
rect 247184 392028 247190 392080
rect 247494 392028 247500 392080
rect 247552 392068 247558 392080
rect 247862 392068 247868 392080
rect 247552 392040 247868 392068
rect 247552 392028 247558 392040
rect 247862 392028 247868 392040
rect 247920 392028 247926 392080
rect 248414 392028 248420 392080
rect 248472 392068 248478 392080
rect 248966 392068 248972 392080
rect 248472 392040 248972 392068
rect 248472 392028 248478 392040
rect 248966 392028 248972 392040
rect 249024 392028 249030 392080
rect 225230 391960 225236 392012
rect 225288 392000 225294 392012
rect 229002 392000 229008 392012
rect 225288 391972 229008 392000
rect 225288 391960 225294 391972
rect 229002 391960 229008 391972
rect 229060 391960 229066 392012
rect 248414 391892 248420 391944
rect 248472 391932 248478 391944
rect 249334 391932 249340 391944
rect 248472 391904 249340 391932
rect 248472 391892 248478 391904
rect 249334 391892 249340 391904
rect 249392 391892 249398 391944
rect 248690 391688 248696 391740
rect 248748 391728 248754 391740
rect 249150 391728 249156 391740
rect 248748 391700 249156 391728
rect 248748 391688 248754 391700
rect 249150 391688 249156 391700
rect 249208 391688 249214 391740
rect 233418 391416 233424 391468
rect 233476 391456 233482 391468
rect 299566 391456 299572 391468
rect 233476 391428 299572 391456
rect 233476 391416 233482 391428
rect 299566 391416 299572 391428
rect 299624 391416 299630 391468
rect 239398 391348 239404 391400
rect 239456 391388 239462 391400
rect 365806 391388 365812 391400
rect 239456 391360 365812 391388
rect 239456 391348 239462 391360
rect 365806 391348 365812 391360
rect 365864 391348 365870 391400
rect 250806 391280 250812 391332
rect 250864 391320 250870 391332
rect 514754 391320 514760 391332
rect 250864 391292 514760 391320
rect 250864 391280 250870 391292
rect 514754 391280 514760 391292
rect 514812 391280 514818 391332
rect 229738 391212 229744 391264
rect 229796 391252 229802 391264
rect 250438 391252 250444 391264
rect 229796 391224 250444 391252
rect 229796 391212 229802 391224
rect 250438 391212 250444 391224
rect 250496 391212 250502 391264
rect 252002 391212 252008 391264
rect 252060 391252 252066 391264
rect 529934 391252 529940 391264
rect 252060 391224 529940 391252
rect 252060 391212 252066 391224
rect 529934 391212 529940 391224
rect 529992 391212 529998 391264
rect 245746 391144 245752 391196
rect 245804 391184 245810 391196
rect 246206 391184 246212 391196
rect 245804 391156 246212 391184
rect 245804 391144 245810 391156
rect 246206 391144 246212 391156
rect 246264 391144 246270 391196
rect 222746 391008 222752 391060
rect 222804 391048 222810 391060
rect 223022 391048 223028 391060
rect 222804 391020 223028 391048
rect 222804 391008 222810 391020
rect 223022 391008 223028 391020
rect 223080 391008 223086 391060
rect 233970 389988 233976 390040
rect 234028 390028 234034 390040
rect 293954 390028 293960 390040
rect 234028 390000 293960 390028
rect 234028 389988 234034 390000
rect 293954 389988 293960 390000
rect 294012 389988 294018 390040
rect 230014 389920 230020 389972
rect 230072 389960 230078 389972
rect 233418 389960 233424 389972
rect 230072 389932 233424 389960
rect 230072 389920 230078 389932
rect 233418 389920 233424 389932
rect 233476 389920 233482 389972
rect 235350 389920 235356 389972
rect 235408 389960 235414 389972
rect 316034 389960 316040 389972
rect 235408 389932 316040 389960
rect 235408 389920 235414 389932
rect 316034 389920 316040 389932
rect 316092 389920 316098 389972
rect 246758 389852 246764 389904
rect 246816 389892 246822 389904
rect 357434 389892 357440 389904
rect 246816 389864 357440 389892
rect 246816 389852 246822 389864
rect 357434 389852 357440 389864
rect 357492 389852 357498 389904
rect 245470 389784 245476 389836
rect 245528 389824 245534 389836
rect 438854 389824 438860 389836
rect 245528 389796 438860 389824
rect 245528 389784 245534 389796
rect 438854 389784 438860 389796
rect 438912 389784 438918 389836
rect 249794 389716 249800 389768
rect 249852 389756 249858 389768
rect 250162 389756 250168 389768
rect 249852 389728 250168 389756
rect 249852 389716 249858 389728
rect 250162 389716 250168 389728
rect 250220 389716 250226 389768
rect 249794 389580 249800 389632
rect 249852 389620 249858 389632
rect 250714 389620 250720 389632
rect 249852 389592 250720 389620
rect 249852 389580 249858 389592
rect 250714 389580 250720 389592
rect 250772 389580 250778 389632
rect 254302 389376 254308 389428
rect 254360 389416 254366 389428
rect 254670 389416 254676 389428
rect 254360 389388 254676 389416
rect 254360 389376 254366 389388
rect 254670 389376 254676 389388
rect 254728 389376 254734 389428
rect 222562 389308 222568 389360
rect 222620 389348 222626 389360
rect 223482 389348 223488 389360
rect 222620 389320 223488 389348
rect 222620 389308 222626 389320
rect 223482 389308 223488 389320
rect 223540 389308 223546 389360
rect 217318 389240 217324 389292
rect 217376 389240 217382 389292
rect 217336 389076 217364 389240
rect 217502 389076 217508 389088
rect 217336 389048 217508 389076
rect 217502 389036 217508 389048
rect 217560 389036 217566 389088
rect 299290 379448 299296 379500
rect 299348 379488 299354 379500
rect 580166 379488 580172 379500
rect 299348 379460 580172 379488
rect 299348 379448 299354 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 98638 372552 98644 372564
rect 3384 372524 98644 372552
rect 3384 372512 3390 372524
rect 98638 372512 98644 372524
rect 98696 372512 98702 372564
rect 296438 365644 296444 365696
rect 296496 365684 296502 365696
rect 580166 365684 580172 365696
rect 296496 365656 580172 365684
rect 296496 365644 296502 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 5166 358476 5172 358488
rect 2832 358448 5172 358476
rect 2832 358436 2838 358448
rect 5166 358436 5172 358448
rect 5224 358436 5230 358488
rect 250346 356804 250352 356856
rect 250404 356844 250410 356856
rect 514846 356844 514852 356856
rect 250404 356816 514852 356844
rect 250404 356804 250410 356816
rect 514846 356804 514852 356816
rect 514904 356804 514910 356856
rect 250530 356736 250536 356788
rect 250588 356776 250594 356788
rect 517514 356776 517520 356788
rect 250588 356748 517520 356776
rect 250588 356736 250594 356748
rect 517514 356736 517520 356748
rect 517572 356736 517578 356788
rect 251818 356668 251824 356720
rect 251876 356708 251882 356720
rect 531314 356708 531320 356720
rect 251876 356680 531320 356708
rect 251876 356668 251882 356680
rect 531314 356668 531320 356680
rect 531372 356668 531378 356720
rect 232590 355580 232596 355632
rect 232648 355620 232654 355632
rect 281534 355620 281540 355632
rect 232648 355592 281540 355620
rect 232648 355580 232654 355592
rect 281534 355580 281540 355592
rect 281592 355580 281598 355632
rect 232498 355512 232504 355564
rect 232556 355552 232562 355564
rect 288434 355552 288440 355564
rect 232556 355524 288440 355552
rect 232556 355512 232562 355524
rect 288434 355512 288440 355524
rect 288492 355512 288498 355564
rect 184934 355444 184940 355496
rect 184992 355484 184998 355496
rect 224218 355484 224224 355496
rect 184992 355456 224224 355484
rect 184992 355444 184998 355456
rect 224218 355444 224224 355456
rect 224276 355444 224282 355496
rect 250162 355444 250168 355496
rect 250220 355484 250226 355496
rect 506474 355484 506480 355496
rect 250220 355456 506480 355484
rect 250220 355444 250226 355456
rect 506474 355444 506480 355456
rect 506532 355444 506538 355496
rect 110414 355376 110420 355428
rect 110472 355416 110478 355428
rect 208026 355416 208032 355428
rect 110472 355388 208032 355416
rect 110472 355376 110478 355388
rect 208026 355376 208032 355388
rect 208084 355376 208090 355428
rect 250254 355376 250260 355428
rect 250312 355416 250318 355428
rect 510614 355416 510620 355428
rect 250312 355388 510620 355416
rect 250312 355376 250318 355388
rect 510614 355376 510620 355388
rect 510672 355376 510678 355428
rect 104894 355308 104900 355360
rect 104952 355348 104958 355360
rect 218514 355348 218520 355360
rect 104952 355320 218520 355348
rect 104952 355308 104958 355320
rect 218514 355308 218520 355320
rect 218572 355308 218578 355360
rect 253290 355308 253296 355360
rect 253348 355348 253354 355360
rect 550634 355348 550640 355360
rect 253348 355320 550640 355348
rect 253348 355308 253354 355320
rect 550634 355308 550640 355320
rect 550692 355308 550698 355360
rect 200114 354560 200120 354612
rect 200172 354600 200178 354612
rect 225414 354600 225420 354612
rect 200172 354572 225420 354600
rect 200172 354560 200178 354572
rect 225414 354560 225420 354572
rect 225472 354560 225478 354612
rect 180794 354492 180800 354544
rect 180852 354532 180858 354544
rect 224126 354532 224132 354544
rect 180852 354504 224132 354532
rect 180852 354492 180858 354504
rect 224126 354492 224132 354504
rect 224184 354492 224190 354544
rect 176654 354424 176660 354476
rect 176712 354464 176718 354476
rect 224034 354464 224040 354476
rect 176712 354436 224040 354464
rect 176712 354424 176718 354436
rect 224034 354424 224040 354436
rect 224092 354424 224098 354476
rect 97994 354356 98000 354408
rect 98052 354396 98058 354408
rect 217134 354396 217140 354408
rect 98052 354368 217140 354396
rect 98052 354356 98058 354368
rect 217134 354356 217140 354368
rect 217192 354356 217198 354408
rect 91094 354288 91100 354340
rect 91152 354328 91158 354340
rect 216950 354328 216956 354340
rect 91152 354300 216956 354328
rect 91152 354288 91158 354300
rect 216950 354288 216956 354300
rect 217008 354288 217014 354340
rect 238110 354288 238116 354340
rect 238168 354328 238174 354340
rect 353294 354328 353300 354340
rect 238168 354300 353300 354328
rect 238168 354288 238174 354300
rect 353294 354288 353300 354300
rect 353352 354288 353358 354340
rect 86954 354220 86960 354272
rect 87012 354260 87018 354272
rect 217042 354260 217048 354272
rect 87012 354232 217048 354260
rect 87012 354220 87018 354232
rect 217042 354220 217048 354232
rect 217100 354220 217106 354272
rect 240870 354220 240876 354272
rect 240928 354260 240934 354272
rect 391934 354260 391940 354272
rect 240928 354232 391940 354260
rect 240928 354220 240934 354232
rect 391934 354220 391940 354232
rect 391992 354220 391998 354272
rect 70394 354152 70400 354204
rect 70452 354192 70458 354204
rect 212074 354192 212080 354204
rect 70452 354164 212080 354192
rect 70452 354152 70458 354164
rect 212074 354152 212080 354164
rect 212132 354152 212138 354204
rect 241974 354152 241980 354204
rect 242032 354192 242038 354204
rect 411254 354192 411260 354204
rect 242032 354164 411260 354192
rect 242032 354152 242038 354164
rect 411254 354152 411260 354164
rect 411312 354152 411318 354204
rect 62114 354084 62120 354136
rect 62172 354124 62178 354136
rect 214558 354124 214564 354136
rect 62172 354096 214564 354124
rect 62172 354084 62178 354096
rect 214558 354084 214564 354096
rect 214616 354084 214622 354136
rect 244826 354084 244832 354136
rect 244884 354124 244890 354136
rect 445754 354124 445760 354136
rect 244884 354096 445760 354124
rect 244884 354084 244890 354096
rect 445754 354084 445760 354096
rect 445812 354084 445818 354136
rect 42794 354016 42800 354068
rect 42852 354056 42858 354068
rect 212994 354056 213000 354068
rect 42852 354028 213000 354056
rect 42852 354016 42858 354028
rect 212994 354016 213000 354028
rect 213052 354016 213058 354068
rect 253198 354016 253204 354068
rect 253256 354056 253262 354068
rect 542354 354056 542360 354068
rect 253256 354028 542360 354056
rect 253256 354016 253262 354028
rect 542354 354016 542360 354028
rect 542412 354016 542418 354068
rect 35894 353948 35900 354000
rect 35952 353988 35958 354000
rect 213086 353988 213092 354000
rect 35952 353960 213092 353988
rect 35952 353948 35958 353960
rect 213086 353948 213092 353960
rect 213144 353948 213150 354000
rect 229646 353948 229652 354000
rect 229704 353988 229710 354000
rect 241790 353988 241796 354000
rect 229704 353960 241796 353988
rect 229704 353948 229710 353960
rect 241790 353948 241796 353960
rect 241848 353948 241854 354000
rect 253106 353948 253112 354000
rect 253164 353988 253170 354000
rect 546494 353988 546500 354000
rect 253164 353960 546500 353988
rect 253164 353948 253170 353960
rect 546494 353948 546500 353960
rect 546552 353948 546558 354000
rect 269850 353200 269856 353252
rect 269908 353240 269914 353252
rect 580166 353240 580172 353252
rect 269908 353212 580172 353240
rect 269908 353200 269914 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 230934 352860 230940 352912
rect 230992 352900 230998 352912
rect 270494 352900 270500 352912
rect 230992 352872 270500 352900
rect 230992 352860 230998 352872
rect 270494 352860 270500 352872
rect 270552 352860 270558 352912
rect 235166 352792 235172 352844
rect 235224 352832 235230 352844
rect 317414 352832 317420 352844
rect 235224 352804 317420 352832
rect 235224 352792 235230 352804
rect 317414 352792 317420 352804
rect 317472 352792 317478 352844
rect 235258 352724 235264 352776
rect 235316 352764 235322 352776
rect 321554 352764 321560 352776
rect 235316 352736 321560 352764
rect 235316 352724 235322 352736
rect 321554 352724 321560 352736
rect 321612 352724 321618 352776
rect 239306 352656 239312 352708
rect 239364 352696 239370 352708
rect 367094 352696 367100 352708
rect 239364 352668 367100 352696
rect 239364 352656 239370 352668
rect 367094 352656 367100 352668
rect 367152 352656 367158 352708
rect 149054 352588 149060 352640
rect 149112 352628 149118 352640
rect 221550 352628 221556 352640
rect 149112 352600 221556 352628
rect 149112 352588 149118 352600
rect 221550 352588 221556 352600
rect 221608 352588 221614 352640
rect 246574 352588 246580 352640
rect 246632 352628 246638 352640
rect 379514 352628 379520 352640
rect 246632 352600 379520 352628
rect 246632 352588 246638 352600
rect 379514 352588 379520 352600
rect 379572 352588 379578 352640
rect 88334 352520 88340 352572
rect 88392 352560 88398 352572
rect 210602 352560 210608 352572
rect 88392 352532 210608 352560
rect 88392 352520 88398 352532
rect 210602 352520 210608 352532
rect 210660 352520 210666 352572
rect 241882 352520 241888 352572
rect 241940 352560 241946 352572
rect 404354 352560 404360 352572
rect 241940 352532 404360 352560
rect 241940 352520 241946 352532
rect 404354 352520 404360 352532
rect 404412 352520 404418 352572
rect 220814 351908 220820 351960
rect 220872 351948 220878 351960
rect 226794 351948 226800 351960
rect 220872 351920 226800 351948
rect 220872 351908 220878 351920
rect 226794 351908 226800 351920
rect 226852 351908 226858 351960
rect 233786 351296 233792 351348
rect 233844 351336 233850 351348
rect 300854 351336 300860 351348
rect 233844 351308 300860 351336
rect 233844 351296 233850 351308
rect 300854 351296 300860 351308
rect 300912 351296 300918 351348
rect 142154 351228 142160 351280
rect 142212 351268 142218 351280
rect 221458 351268 221464 351280
rect 142212 351240 221464 351268
rect 142212 351228 142218 351240
rect 221458 351228 221464 351240
rect 221516 351228 221522 351280
rect 242618 351228 242624 351280
rect 242676 351268 242682 351280
rect 393314 351268 393320 351280
rect 242676 351240 393320 351268
rect 242676 351228 242682 351240
rect 393314 351228 393320 351240
rect 393372 351228 393378 351280
rect 74534 351160 74540 351212
rect 74592 351200 74598 351212
rect 216122 351200 216128 351212
rect 74592 351172 216128 351200
rect 74592 351160 74598 351172
rect 216122 351160 216128 351172
rect 216180 351160 216186 351212
rect 218514 351160 218520 351212
rect 218572 351200 218578 351212
rect 226702 351200 226708 351212
rect 218572 351172 226708 351200
rect 218572 351160 218578 351172
rect 226702 351160 226708 351172
rect 226760 351160 226766 351212
rect 243630 351160 243636 351212
rect 243688 351200 243694 351212
rect 423674 351200 423680 351212
rect 243688 351172 423680 351200
rect 243688 351160 243694 351172
rect 423674 351160 423680 351172
rect 423732 351160 423738 351212
rect 254486 348372 254492 348424
rect 254544 348412 254550 348424
rect 572714 348412 572720 348424
rect 254544 348384 572720 348412
rect 254544 348372 254550 348384
rect 572714 348372 572720 348384
rect 572772 348372 572778 348424
rect 23474 338716 23480 338768
rect 23532 338756 23538 338768
rect 209222 338756 209228 338768
rect 23532 338728 209228 338756
rect 23532 338716 23538 338728
rect 209222 338716 209228 338728
rect 209280 338716 209286 338768
rect 260098 335996 260104 336048
rect 260156 336036 260162 336048
rect 449894 336036 449900 336048
rect 260156 336008 449900 336036
rect 260156 335996 260162 336008
rect 449894 335996 449900 336008
rect 449952 335996 449958 336048
rect 257614 334568 257620 334620
rect 257672 334608 257678 334620
rect 429194 334608 429200 334620
rect 257672 334580 429200 334608
rect 257672 334568 257678 334580
rect 429194 334568 429200 334580
rect 429252 334568 429258 334620
rect 299106 325592 299112 325644
rect 299164 325632 299170 325644
rect 580166 325632 580172 325644
rect 299164 325604 580172 325632
rect 299164 325592 299170 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 199654 320124 199660 320136
rect 3384 320096 199660 320124
rect 3384 320084 3390 320096
rect 199654 320084 199660 320096
rect 199712 320084 199718 320136
rect 296254 313216 296260 313268
rect 296312 313256 296318 313268
rect 580166 313256 580172 313268
rect 296312 313228 580172 313256
rect 296312 313216 296318 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 2774 306212 2780 306264
rect 2832 306252 2838 306264
rect 5074 306252 5080 306264
rect 2832 306224 5080 306252
rect 2832 306212 2838 306224
rect 5074 306212 5080 306224
rect 5132 306212 5138 306264
rect 258810 305600 258816 305652
rect 258868 305640 258874 305652
rect 436094 305640 436100 305652
rect 258868 305612 436100 305640
rect 258868 305600 258874 305612
rect 436094 305600 436100 305612
rect 436152 305600 436158 305652
rect 265986 299412 265992 299464
rect 266044 299452 266050 299464
rect 580166 299452 580172 299464
rect 266044 299424 580172 299452
rect 266044 299412 266050 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 299198 273164 299204 273216
rect 299256 273204 299262 273216
rect 580166 273204 580172 273216
rect 299256 273176 580172 273204
rect 299256 273164 299262 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3142 267656 3148 267708
rect 3200 267696 3206 267708
rect 196710 267696 196716 267708
rect 3200 267668 196716 267696
rect 3200 267656 3206 267668
rect 196710 267656 196716 267668
rect 196768 267656 196774 267708
rect 296346 259360 296352 259412
rect 296404 259400 296410 259412
rect 580166 259400 580172 259412
rect 296404 259372 580172 259400
rect 296404 259360 296410 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 268378 245556 268384 245608
rect 268436 245596 268442 245608
rect 580166 245596 580172 245608
rect 268436 245568 580172 245596
rect 268436 245556 268442 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 298922 233180 298928 233232
rect 298980 233220 298986 233232
rect 579982 233220 579988 233232
rect 298980 233192 579988 233220
rect 298980 233180 298986 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 296162 219376 296168 219428
rect 296220 219416 296226 219428
rect 580166 219416 580172 219428
rect 296220 219388 580172 219416
rect 296220 219376 296226 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3050 215228 3056 215280
rect 3108 215268 3114 215280
rect 199562 215268 199568 215280
rect 3108 215240 199568 215268
rect 3108 215228 3114 215240
rect 199562 215228 199568 215240
rect 199620 215228 199626 215280
rect 299014 206932 299020 206984
rect 299072 206972 299078 206984
rect 579798 206972 579804 206984
rect 299072 206944 579804 206972
rect 299072 206932 299078 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 2774 202648 2780 202700
rect 2832 202688 2838 202700
rect 4982 202688 4988 202700
rect 2832 202660 4988 202688
rect 2832 202648 2838 202660
rect 4982 202648 4988 202660
rect 5040 202648 5046 202700
rect 298830 193128 298836 193180
rect 298888 193168 298894 193180
rect 580166 193168 580172 193180
rect 298888 193140 580172 193168
rect 298888 193128 298894 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 275370 191088 275376 191140
rect 275428 191128 275434 191140
rect 582374 191128 582380 191140
rect 275428 191100 582380 191128
rect 275428 191088 275434 191100
rect 582374 191088 582380 191100
rect 582432 191088 582438 191140
rect 264330 188300 264336 188352
rect 264388 188340 264394 188352
rect 460934 188340 460940 188352
rect 264388 188312 460940 188340
rect 264388 188300 264394 188312
rect 460934 188300 460940 188312
rect 460992 188300 460998 188352
rect 261478 186940 261484 186992
rect 261536 186980 261542 186992
rect 442994 186980 443000 186992
rect 261536 186952 443000 186980
rect 261536 186940 261542 186952
rect 442994 186940 443000 186952
rect 443052 186940 443058 186992
rect 38654 180072 38660 180124
rect 38712 180112 38718 180124
rect 202138 180112 202144 180124
rect 38712 180084 202144 180112
rect 38712 180072 38718 180084
rect 202138 180072 202144 180084
rect 202196 180072 202202 180124
rect 295978 179324 295984 179376
rect 296036 179364 296042 179376
rect 580166 179364 580172 179376
rect 296036 179336 580172 179364
rect 296036 179324 296042 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 102226 178644 102232 178696
rect 102284 178684 102290 178696
rect 207934 178684 207940 178696
rect 102284 178656 207940 178684
rect 102284 178644 102290 178656
rect 207934 178644 207940 178656
rect 207992 178644 207998 178696
rect 240778 178644 240784 178696
rect 240836 178684 240842 178696
rect 389174 178684 389180 178696
rect 240836 178656 389180 178684
rect 240836 178644 240842 178656
rect 389174 178644 389180 178656
rect 389232 178644 389238 178696
rect 155954 177556 155960 177608
rect 156012 177596 156018 177608
rect 222930 177596 222936 177608
rect 156012 177568 222936 177596
rect 156012 177556 156018 177568
rect 222930 177556 222936 177568
rect 222988 177556 222994 177608
rect 124214 177488 124220 177540
rect 124272 177528 124278 177540
rect 219986 177528 219992 177540
rect 124272 177500 219992 177528
rect 124272 177488 124278 177500
rect 219986 177488 219992 177500
rect 220044 177488 220050 177540
rect 111794 177420 111800 177472
rect 111852 177460 111858 177472
rect 218606 177460 218612 177472
rect 111852 177432 218612 177460
rect 111852 177420 111858 177432
rect 218606 177420 218612 177432
rect 218664 177420 218670 177472
rect 80054 177352 80060 177404
rect 80112 177392 80118 177404
rect 216030 177392 216036 177404
rect 80112 177364 216036 177392
rect 80112 177352 80118 177364
rect 216030 177352 216036 177364
rect 216088 177352 216094 177404
rect 228266 177352 228272 177404
rect 228324 177392 228330 177404
rect 232498 177392 232504 177404
rect 228324 177364 232504 177392
rect 228324 177352 228330 177364
rect 232498 177352 232504 177364
rect 232556 177352 232562 177404
rect 9674 177284 9680 177336
rect 9732 177324 9738 177336
rect 210326 177324 210332 177336
rect 9732 177296 210332 177324
rect 9732 177284 9738 177296
rect 210326 177284 210332 177296
rect 210384 177284 210390 177336
rect 228358 177284 228364 177336
rect 228416 177324 228422 177336
rect 235166 177324 235172 177336
rect 228416 177296 235172 177324
rect 228416 177284 228422 177296
rect 235166 177284 235172 177296
rect 235224 177284 235230 177336
rect 242250 177284 242256 177336
rect 242308 177324 242314 177336
rect 372614 177324 372620 177336
rect 242308 177296 372620 177324
rect 242308 177284 242314 177296
rect 372614 177284 372620 177296
rect 372672 177284 372678 177336
rect 31754 168988 31760 169040
rect 31812 169028 31818 169040
rect 203610 169028 203616 169040
rect 31812 169000 203616 169028
rect 31812 168988 31818 169000
rect 203610 168988 203616 169000
rect 203668 168988 203674 169040
rect 269758 167628 269764 167680
rect 269816 167668 269822 167680
rect 581086 167668 581092 167680
rect 269816 167640 581092 167668
rect 269816 167628 269822 167640
rect 581086 167628 581092 167640
rect 581144 167628 581150 167680
rect 275278 166948 275284 167000
rect 275336 166988 275342 167000
rect 580166 166988 580172 167000
rect 275336 166960 580172 166988
rect 275336 166948 275342 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3050 164160 3056 164212
rect 3108 164200 3114 164212
rect 196618 164200 196624 164212
rect 3108 164172 196624 164200
rect 3108 164160 3114 164172
rect 196618 164160 196624 164172
rect 196676 164160 196682 164212
rect 278038 153144 278044 153196
rect 278096 153184 278102 153196
rect 580166 153184 580172 153196
rect 278096 153156 580172 153184
rect 278096 153144 278102 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 2774 149880 2780 149932
rect 2832 149920 2838 149932
rect 4890 149920 4896 149932
rect 2832 149892 4896 149920
rect 2832 149880 2838 149892
rect 4890 149880 4896 149892
rect 4948 149880 4954 149932
rect 265894 139340 265900 139392
rect 265952 139380 265958 139392
rect 580166 139380 580172 139392
rect 265952 139352 580172 139380
rect 265952 139340 265958 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 273898 126896 273904 126948
rect 273956 126936 273962 126948
rect 580166 126936 580172 126948
rect 273956 126908 580172 126936
rect 273956 126896 273962 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 298738 113092 298744 113144
rect 298796 113132 298802 113144
rect 579798 113132 579804 113144
rect 298796 113104 579804 113132
rect 298796 113092 298802 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 199470 111772 199476 111784
rect 3384 111744 199476 111772
rect 3384 111732 3390 111744
rect 199470 111732 199476 111744
rect 199528 111732 199534 111784
rect 296070 100648 296076 100700
rect 296128 100688 296134 100700
rect 580166 100688 580172 100700
rect 296128 100660 580172 100688
rect 296128 100648 296134 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 216950 88952 216956 89004
rect 217008 88992 217014 89004
rect 224954 88992 224960 89004
rect 217008 88964 224960 88992
rect 217008 88952 217014 88964
rect 224954 88952 224960 88964
rect 225012 88952 225018 89004
rect 232406 87728 232412 87780
rect 232464 87768 232470 87780
rect 287054 87768 287060 87780
rect 232464 87740 287060 87768
rect 232464 87728 232470 87740
rect 287054 87728 287060 87740
rect 287112 87728 287118 87780
rect 243538 87660 243544 87712
rect 243596 87700 243602 87712
rect 427814 87700 427820 87712
rect 243596 87672 427820 87700
rect 243596 87660 243602 87672
rect 427814 87660 427820 87672
rect 427872 87660 427878 87712
rect 251726 87592 251732 87644
rect 251784 87632 251790 87644
rect 531406 87632 531412 87644
rect 251784 87604 531412 87632
rect 251784 87592 251790 87604
rect 531406 87592 531412 87604
rect 531464 87592 531470 87644
rect 265802 86912 265808 86964
rect 265860 86952 265866 86964
rect 580166 86952 580172 86964
rect 265860 86924 580172 86952
rect 265860 86912 265866 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 240686 86300 240692 86352
rect 240744 86340 240750 86352
rect 385034 86340 385040 86352
rect 240744 86312 385040 86340
rect 240744 86300 240750 86312
rect 385034 86300 385040 86312
rect 385092 86300 385098 86352
rect 117314 86232 117320 86284
rect 117372 86272 117378 86284
rect 206278 86272 206284 86284
rect 117372 86244 206284 86272
rect 117372 86232 117378 86244
rect 206278 86232 206284 86244
rect 206336 86232 206342 86284
rect 246206 86232 246212 86284
rect 246264 86272 246270 86284
rect 454034 86272 454040 86284
rect 246264 86244 454040 86272
rect 246264 86232 246270 86244
rect 454034 86232 454040 86244
rect 454092 86232 454098 86284
rect 238018 84804 238024 84856
rect 238076 84844 238082 84856
rect 354674 84844 354680 84856
rect 238076 84816 354680 84844
rect 238076 84804 238082 84816
rect 354674 84804 354680 84816
rect 354732 84804 354738 84856
rect 233694 83580 233700 83632
rect 233752 83620 233758 83632
rect 298094 83620 298100 83632
rect 233752 83592 298100 83620
rect 233752 83580 233758 83592
rect 298094 83580 298100 83592
rect 298152 83580 298158 83632
rect 256602 83512 256608 83564
rect 256660 83552 256666 83564
rect 422294 83552 422300 83564
rect 256660 83524 422300 83552
rect 256660 83512 256666 83524
rect 422294 83512 422300 83524
rect 422352 83512 422358 83564
rect 243446 83444 243452 83496
rect 243504 83484 243510 83496
rect 420914 83484 420920 83496
rect 243504 83456 420920 83484
rect 243504 83444 243510 83456
rect 420914 83444 420920 83456
rect 420972 83444 420978 83496
rect 95234 82084 95240 82136
rect 95292 82124 95298 82136
rect 207842 82124 207848 82136
rect 95292 82096 207848 82124
rect 95292 82084 95298 82096
rect 207842 82084 207848 82096
rect 207900 82084 207906 82136
rect 249058 82084 249064 82136
rect 249116 82124 249122 82136
rect 499574 82124 499580 82136
rect 249116 82096 499580 82124
rect 249116 82084 249122 82096
rect 499574 82084 499580 82096
rect 499632 82084 499638 82136
rect 236546 80656 236552 80708
rect 236604 80696 236610 80708
rect 336734 80696 336740 80708
rect 236604 80668 336740 80696
rect 236604 80656 236610 80668
rect 336734 80656 336740 80668
rect 336792 80656 336798 80708
rect 265710 73108 265716 73160
rect 265768 73148 265774 73160
rect 580166 73148 580172 73160
rect 265768 73120 580172 73148
rect 265768 73108 265774 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 257522 71720 257528 71732
rect 3384 71692 257528 71720
rect 3384 71680 3390 71692
rect 257522 71680 257528 71692
rect 257580 71680 257586 71732
rect 283558 60664 283564 60716
rect 283616 60704 283622 60716
rect 580166 60704 580172 60716
rect 283616 60676 580172 60704
rect 283616 60664 283622 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 265618 46860 265624 46912
rect 265676 46900 265682 46912
rect 580166 46900 580172 46912
rect 265676 46872 580172 46900
rect 265676 46860 265682 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 162854 46248 162860 46300
rect 162912 46288 162918 46300
rect 222746 46288 222752 46300
rect 162912 46260 222752 46288
rect 162912 46248 162918 46260
rect 222746 46248 222752 46260
rect 222804 46248 222810 46300
rect 146294 46180 146300 46232
rect 146352 46220 146358 46232
rect 221366 46220 221372 46232
rect 146352 46192 221372 46220
rect 146352 46180 146358 46192
rect 221366 46180 221372 46192
rect 221424 46180 221430 46232
rect 229554 46180 229560 46232
rect 229612 46220 229618 46232
rect 249058 46220 249064 46232
rect 229612 46192 249064 46220
rect 229612 46180 229618 46192
rect 249058 46180 249064 46192
rect 249116 46180 249122 46232
rect 271138 31016 271144 31068
rect 271196 31056 271202 31068
rect 474734 31056 474740 31068
rect 271196 31028 474740 31056
rect 271196 31016 271202 31028
rect 474734 31016 474740 31028
rect 474792 31016 474798 31068
rect 264238 29588 264244 29640
rect 264296 29628 264302 29640
rect 456794 29628 456800 29640
rect 264296 29600 456800 29628
rect 264296 29588 264302 29600
rect 456794 29588 456800 29600
rect 456852 29588 456858 29640
rect 256510 27072 256516 27124
rect 256568 27112 256574 27124
rect 400214 27112 400220 27124
rect 256568 27084 400220 27112
rect 256568 27072 256574 27084
rect 400214 27072 400220 27084
rect 400272 27072 400278 27124
rect 256418 27004 256424 27056
rect 256476 27044 256482 27056
rect 407114 27044 407120 27056
rect 256476 27016 407120 27044
rect 256476 27004 256482 27016
rect 407114 27004 407120 27016
rect 407172 27004 407178 27056
rect 244734 26936 244740 26988
rect 244792 26976 244798 26988
rect 447134 26976 447140 26988
rect 244792 26948 447140 26976
rect 244792 26936 244798 26948
rect 447134 26936 447140 26948
rect 447192 26936 447198 26988
rect 247586 26868 247592 26920
rect 247644 26908 247650 26920
rect 471974 26908 471980 26920
rect 247644 26880 471980 26908
rect 247644 26868 247650 26880
rect 471974 26868 471980 26880
rect 472032 26868 472038 26920
rect 232314 25916 232320 25968
rect 232372 25956 232378 25968
rect 280154 25956 280160 25968
rect 232372 25928 280160 25956
rect 232372 25916 232378 25928
rect 280154 25916 280160 25928
rect 280212 25916 280218 25968
rect 232222 25848 232228 25900
rect 232280 25888 232286 25900
rect 284294 25888 284300 25900
rect 232280 25860 284300 25888
rect 232280 25848 232286 25860
rect 284294 25848 284300 25860
rect 284352 25848 284358 25900
rect 235074 25780 235080 25832
rect 235132 25820 235138 25832
rect 311894 25820 311900 25832
rect 235132 25792 311900 25820
rect 235132 25780 235138 25792
rect 311894 25780 311900 25792
rect 311952 25780 311958 25832
rect 234982 25712 234988 25764
rect 235040 25752 235046 25764
rect 318794 25752 318800 25764
rect 235040 25724 318800 25752
rect 235040 25712 235046 25724
rect 318794 25712 318800 25724
rect 318852 25712 318858 25764
rect 240594 25644 240600 25696
rect 240652 25684 240658 25696
rect 390554 25684 390560 25696
rect 240652 25656 390560 25684
rect 240652 25644 240658 25656
rect 390554 25644 390560 25656
rect 390612 25644 390618 25696
rect 243354 25576 243360 25628
rect 243412 25616 243418 25628
rect 425054 25616 425060 25628
rect 243412 25588 425060 25616
rect 243412 25576 243418 25588
rect 425054 25576 425060 25588
rect 425112 25576 425118 25628
rect 254394 25508 254400 25560
rect 254452 25548 254458 25560
rect 567194 25548 567200 25560
rect 254452 25520 567200 25548
rect 254452 25508 254458 25520
rect 567194 25508 567200 25520
rect 567252 25508 567258 25560
rect 246114 24420 246120 24472
rect 246172 24460 246178 24472
rect 463694 24460 463700 24472
rect 246172 24432 463700 24460
rect 246172 24420 246178 24432
rect 463694 24420 463700 24432
rect 463752 24420 463758 24472
rect 247310 24352 247316 24404
rect 247368 24392 247374 24404
rect 473354 24392 473360 24404
rect 247368 24364 473360 24392
rect 247368 24352 247374 24364
rect 473354 24352 473360 24364
rect 473412 24352 473418 24404
rect 247402 24284 247408 24336
rect 247460 24324 247466 24336
rect 477494 24324 477500 24336
rect 247460 24296 477500 24324
rect 247460 24284 247466 24296
rect 477494 24284 477500 24296
rect 477552 24284 477558 24336
rect 247494 24216 247500 24268
rect 247552 24256 247558 24268
rect 481634 24256 481640 24268
rect 247552 24228 481640 24256
rect 247552 24216 247558 24228
rect 481634 24216 481640 24228
rect 481692 24216 481698 24268
rect 248966 24148 248972 24200
rect 249024 24188 249030 24200
rect 490006 24188 490012 24200
rect 249024 24160 490012 24188
rect 249024 24148 249030 24160
rect 490006 24148 490012 24160
rect 490064 24148 490070 24200
rect 248874 24080 248880 24132
rect 248932 24120 248938 24132
rect 496814 24120 496820 24132
rect 248932 24092 496820 24120
rect 248932 24080 248938 24092
rect 496814 24080 496820 24092
rect 496872 24080 496878 24132
rect 244918 23060 244924 23112
rect 244976 23100 244982 23112
rect 386414 23100 386420 23112
rect 244976 23072 386420 23100
rect 244976 23060 244982 23072
rect 386414 23060 386420 23072
rect 386472 23060 386478 23112
rect 241698 22992 241704 23044
rect 241756 23032 241762 23044
rect 407206 23032 407212 23044
rect 241756 23004 407212 23032
rect 241756 22992 241762 23004
rect 407206 22992 407212 23004
rect 407264 22992 407270 23044
rect 244550 22924 244556 22976
rect 244608 22964 244614 22976
rect 441614 22964 441620 22976
rect 244608 22936 441620 22964
rect 244608 22924 244614 22936
rect 441614 22924 441620 22936
rect 441672 22924 441678 22976
rect 244642 22856 244648 22908
rect 244700 22896 244706 22908
rect 448514 22896 448520 22908
rect 244700 22868 448520 22896
rect 244700 22856 244706 22868
rect 448514 22856 448520 22868
rect 448572 22856 448578 22908
rect 245930 22788 245936 22840
rect 245988 22828 245994 22840
rect 456886 22828 456892 22840
rect 245988 22800 456892 22828
rect 245988 22788 245994 22800
rect 456886 22788 456892 22800
rect 456944 22788 456950 22840
rect 246022 22720 246028 22772
rect 246080 22760 246086 22772
rect 459554 22760 459560 22772
rect 246080 22732 459560 22760
rect 246080 22720 246086 22732
rect 459554 22720 459560 22732
rect 459612 22720 459618 22772
rect 236454 21700 236460 21752
rect 236512 21740 236518 21752
rect 335354 21740 335360 21752
rect 236512 21712 335360 21740
rect 236512 21700 236518 21712
rect 335354 21700 335360 21712
rect 335412 21700 335418 21752
rect 236362 21632 236368 21684
rect 236420 21672 236426 21684
rect 339494 21672 339500 21684
rect 236420 21644 339500 21672
rect 236420 21632 236426 21644
rect 339494 21632 339500 21644
rect 339552 21632 339558 21684
rect 237926 21564 237932 21616
rect 237984 21604 237990 21616
rect 349154 21604 349160 21616
rect 237984 21576 349160 21604
rect 237984 21564 237990 21576
rect 349154 21564 349160 21576
rect 349212 21564 349218 21616
rect 237834 21496 237840 21548
rect 237892 21536 237898 21548
rect 357526 21536 357532 21548
rect 237892 21508 357532 21536
rect 237892 21496 237898 21508
rect 357526 21496 357532 21508
rect 357584 21496 357590 21548
rect 239214 21428 239220 21480
rect 239272 21468 239278 21480
rect 371234 21468 371240 21480
rect 239272 21440 371240 21468
rect 239272 21428 239278 21440
rect 371234 21428 371240 21440
rect 371292 21428 371298 21480
rect 239122 21360 239128 21412
rect 239180 21400 239186 21412
rect 373994 21400 374000 21412
rect 239180 21372 374000 21400
rect 239180 21360 239186 21372
rect 373994 21360 374000 21372
rect 374052 21360 374058 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 199378 20652 199384 20664
rect 3476 20624 199384 20652
rect 3476 20612 3482 20624
rect 199378 20612 199384 20624
rect 199436 20612 199442 20664
rect 232130 20204 232136 20256
rect 232188 20244 232194 20256
rect 285674 20244 285680 20256
rect 232188 20216 285680 20244
rect 232188 20204 232194 20216
rect 285674 20204 285680 20216
rect 285732 20204 285738 20256
rect 233602 20136 233608 20188
rect 233660 20176 233666 20188
rect 296714 20176 296720 20188
rect 233660 20148 296720 20176
rect 233660 20136 233666 20148
rect 296714 20136 296720 20148
rect 296772 20136 296778 20188
rect 234890 20068 234896 20120
rect 234948 20108 234954 20120
rect 314654 20108 314660 20120
rect 234948 20080 314660 20108
rect 234948 20068 234954 20080
rect 314654 20068 314660 20080
rect 314712 20068 314718 20120
rect 236270 20000 236276 20052
rect 236328 20040 236334 20052
rect 332686 20040 332692 20052
rect 236328 20012 332692 20040
rect 236328 20000 236334 20012
rect 332686 20000 332692 20012
rect 332744 20000 332750 20052
rect 255406 19932 255412 19984
rect 255464 19972 255470 19984
rect 578234 19972 578240 19984
rect 255464 19944 578240 19972
rect 255464 19932 255470 19944
rect 578234 19932 578240 19944
rect 578292 19932 578298 19984
rect 230842 19116 230848 19168
rect 230900 19156 230906 19168
rect 267826 19156 267832 19168
rect 230900 19128 267832 19156
rect 230900 19116 230906 19128
rect 267826 19116 267832 19128
rect 267884 19116 267890 19168
rect 233878 19048 233884 19100
rect 233936 19088 233942 19100
rect 271874 19088 271880 19100
rect 233936 19060 271880 19088
rect 233936 19048 233942 19060
rect 271874 19048 271880 19060
rect 271932 19048 271938 19100
rect 232038 18980 232044 19032
rect 232096 19020 232102 19032
rect 278774 19020 278780 19032
rect 232096 18992 278780 19020
rect 232096 18980 232102 18992
rect 278774 18980 278780 18992
rect 278832 18980 278838 19032
rect 231946 18912 231952 18964
rect 232004 18952 232010 18964
rect 282914 18952 282920 18964
rect 232004 18924 282920 18952
rect 232004 18912 232010 18924
rect 282914 18912 282920 18924
rect 282972 18912 282978 18964
rect 233510 18844 233516 18896
rect 233568 18884 233574 18896
rect 303614 18884 303620 18896
rect 233568 18856 303620 18884
rect 233568 18844 233574 18856
rect 303614 18844 303620 18856
rect 303672 18844 303678 18896
rect 240502 18776 240508 18828
rect 240560 18816 240566 18828
rect 396074 18816 396080 18828
rect 240560 18788 396080 18816
rect 240560 18776 240566 18788
rect 396074 18776 396080 18788
rect 396132 18776 396138 18828
rect 243262 18708 243268 18760
rect 243320 18748 243326 18760
rect 418154 18748 418160 18760
rect 243320 18720 418160 18748
rect 243320 18708 243326 18720
rect 418154 18708 418160 18720
rect 418212 18708 418218 18760
rect 254210 18640 254216 18692
rect 254268 18680 254274 18692
rect 563054 18680 563060 18692
rect 254268 18652 563060 18680
rect 254268 18640 254274 18652
rect 563054 18640 563060 18652
rect 563112 18640 563118 18692
rect 254302 18572 254308 18624
rect 254360 18612 254366 18624
rect 569954 18612 569960 18624
rect 254360 18584 569960 18612
rect 254360 18572 254366 18584
rect 569954 18572 569960 18584
rect 570012 18572 570018 18624
rect 240410 17552 240416 17604
rect 240468 17592 240474 17604
rect 397454 17592 397460 17604
rect 240468 17564 397460 17592
rect 240468 17552 240474 17564
rect 397454 17552 397460 17564
rect 397512 17552 397518 17604
rect 251542 17484 251548 17536
rect 251600 17524 251606 17536
rect 527174 17524 527180 17536
rect 251600 17496 527180 17524
rect 251600 17484 251606 17496
rect 527174 17484 527180 17496
rect 527232 17484 527238 17536
rect 251634 17416 251640 17468
rect 251692 17456 251698 17468
rect 534074 17456 534080 17468
rect 251692 17428 534080 17456
rect 251692 17416 251698 17428
rect 534074 17416 534080 17428
rect 534132 17416 534138 17468
rect 253014 17348 253020 17400
rect 253072 17388 253078 17400
rect 545114 17388 545120 17400
rect 253072 17360 545120 17388
rect 253072 17348 253078 17360
rect 545114 17348 545120 17360
rect 545172 17348 545178 17400
rect 252830 17280 252836 17332
rect 252888 17320 252894 17332
rect 547874 17320 547880 17332
rect 252888 17292 547880 17320
rect 252888 17280 252894 17292
rect 547874 17280 547880 17292
rect 547932 17280 547938 17332
rect 252922 17212 252928 17264
rect 252980 17252 252986 17264
rect 552014 17252 552020 17264
rect 252980 17224 552020 17252
rect 252980 17212 252986 17224
rect 552014 17212 552020 17224
rect 552072 17212 552078 17264
rect 239030 16260 239036 16312
rect 239088 16300 239094 16312
rect 376018 16300 376024 16312
rect 239088 16272 376024 16300
rect 239088 16260 239094 16272
rect 376018 16260 376024 16272
rect 376076 16260 376082 16312
rect 248598 16192 248604 16244
rect 248656 16232 248662 16244
rect 495434 16232 495440 16244
rect 248656 16204 495440 16232
rect 248656 16192 248662 16204
rect 495434 16192 495440 16204
rect 495492 16192 495498 16244
rect 198734 16124 198740 16176
rect 198792 16164 198798 16176
rect 225322 16164 225328 16176
rect 198792 16136 225328 16164
rect 198792 16124 198798 16136
rect 225322 16124 225328 16136
rect 225380 16124 225386 16176
rect 248690 16124 248696 16176
rect 248748 16164 248754 16176
rect 498930 16164 498936 16176
rect 248748 16136 498936 16164
rect 248748 16124 248754 16136
rect 498930 16124 498936 16136
rect 498988 16124 498994 16176
rect 123018 16056 123024 16108
rect 123076 16096 123082 16108
rect 219894 16096 219900 16108
rect 123076 16068 219900 16096
rect 123076 16056 123082 16068
rect 219894 16056 219900 16068
rect 219952 16056 219958 16108
rect 248782 16056 248788 16108
rect 248840 16096 248846 16108
rect 502978 16096 502984 16108
rect 248840 16068 502984 16096
rect 248840 16056 248846 16068
rect 502978 16056 502984 16068
rect 503036 16056 503042 16108
rect 114002 15988 114008 16040
rect 114060 16028 114066 16040
rect 218422 16028 218428 16040
rect 114060 16000 218428 16028
rect 114060 15988 114066 16000
rect 218422 15988 218428 16000
rect 218480 15988 218486 16040
rect 249886 15988 249892 16040
rect 249944 16028 249950 16040
rect 509602 16028 509608 16040
rect 249944 16000 509608 16028
rect 249944 15988 249950 16000
rect 509602 15988 509608 16000
rect 509660 15988 509666 16040
rect 85666 15920 85672 15972
rect 85724 15960 85730 15972
rect 210510 15960 210516 15972
rect 85724 15932 210516 15960
rect 85724 15920 85730 15932
rect 210510 15920 210516 15932
rect 210568 15920 210574 15972
rect 250070 15920 250076 15972
rect 250128 15960 250134 15972
rect 513374 15960 513380 15972
rect 250128 15932 513380 15960
rect 250128 15920 250134 15932
rect 513374 15920 513380 15932
rect 513432 15920 513438 15972
rect 60826 15852 60832 15904
rect 60884 15892 60890 15904
rect 211890 15892 211896 15904
rect 60884 15864 211896 15892
rect 60884 15852 60890 15864
rect 211890 15852 211896 15864
rect 211948 15852 211954 15904
rect 249978 15852 249984 15904
rect 250036 15892 250042 15904
rect 517146 15892 517152 15904
rect 250036 15864 517152 15892
rect 250036 15852 250042 15864
rect 517146 15852 517152 15864
rect 517204 15852 517210 15904
rect 56778 14832 56784 14884
rect 56836 14872 56842 14884
rect 214466 14872 214472 14884
rect 56836 14844 214472 14872
rect 56836 14832 56842 14844
rect 214466 14832 214472 14844
rect 214524 14832 214530 14884
rect 45002 14764 45008 14816
rect 45060 14804 45066 14816
rect 212810 14804 212816 14816
rect 45060 14776 212816 14804
rect 45060 14764 45066 14776
rect 212810 14764 212816 14776
rect 212868 14764 212874 14816
rect 238938 14764 238944 14816
rect 238996 14804 239002 14816
rect 369394 14804 369400 14816
rect 238996 14776 369400 14804
rect 238996 14764 239002 14776
rect 369394 14764 369400 14776
rect 369452 14764 369458 14816
rect 41874 14696 41880 14748
rect 41932 14736 41938 14748
rect 211154 14736 211160 14748
rect 41932 14708 211160 14736
rect 41932 14696 41938 14708
rect 211154 14696 211160 14708
rect 211212 14696 211218 14748
rect 246942 14696 246948 14748
rect 247000 14736 247006 14748
rect 462314 14736 462320 14748
rect 247000 14708 462320 14736
rect 247000 14696 247006 14708
rect 462314 14696 462320 14708
rect 462372 14696 462378 14748
rect 38378 14628 38384 14680
rect 38436 14668 38442 14680
rect 212902 14668 212908 14680
rect 38436 14640 212908 14668
rect 38436 14628 38442 14640
rect 212902 14628 212908 14640
rect 212960 14628 212966 14680
rect 245838 14628 245844 14680
rect 245896 14668 245902 14680
rect 465810 14668 465816 14680
rect 245896 14640 465816 14668
rect 245896 14628 245902 14640
rect 465810 14628 465816 14640
rect 465868 14628 465874 14680
rect 34514 14560 34520 14612
rect 34572 14600 34578 14612
rect 211798 14600 211804 14612
rect 34572 14572 211804 14600
rect 34572 14560 34578 14572
rect 211798 14560 211804 14572
rect 211856 14560 211862 14612
rect 247034 14560 247040 14612
rect 247092 14600 247098 14612
rect 473446 14600 473452 14612
rect 247092 14572 473452 14600
rect 247092 14560 247098 14572
rect 473446 14560 473452 14572
rect 473504 14560 473510 14612
rect 22554 14492 22560 14544
rect 22612 14532 22618 14544
rect 211338 14532 211344 14544
rect 22612 14504 211344 14532
rect 22612 14492 22618 14504
rect 211338 14492 211344 14504
rect 211396 14492 211402 14544
rect 247218 14492 247224 14544
rect 247276 14532 247282 14544
rect 476482 14532 476488 14544
rect 247276 14504 476488 14532
rect 247276 14492 247282 14504
rect 476482 14492 476488 14504
rect 476540 14492 476546 14544
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 211430 14464 211436 14476
rect 18012 14436 211436 14464
rect 18012 14424 18018 14436
rect 211430 14424 211436 14436
rect 211488 14424 211494 14476
rect 247126 14424 247132 14476
rect 247184 14464 247190 14476
rect 481726 14464 481732 14476
rect 247184 14436 481732 14464
rect 247184 14424 247190 14436
rect 481726 14424 481732 14436
rect 481784 14424 481790 14476
rect 133138 13540 133144 13592
rect 133196 13580 133202 13592
rect 215662 13580 215668 13592
rect 133196 13552 215668 13580
rect 133196 13540 133202 13552
rect 215662 13540 215668 13552
rect 215720 13540 215726 13592
rect 73338 13472 73344 13524
rect 73396 13512 73402 13524
rect 215754 13512 215760 13524
rect 73396 13484 215760 13512
rect 73396 13472 73402 13484
rect 215754 13472 215760 13484
rect 215812 13472 215818 13524
rect 69842 13404 69848 13456
rect 69900 13444 69906 13456
rect 215846 13444 215852 13456
rect 69900 13416 215852 13444
rect 69900 13404 69906 13416
rect 215846 13404 215852 13416
rect 215904 13404 215910 13456
rect 237742 13404 237748 13456
rect 237800 13444 237806 13456
rect 351178 13444 351184 13456
rect 237800 13416 351184 13444
rect 237800 13404 237806 13416
rect 351178 13404 351184 13416
rect 351236 13404 351242 13456
rect 59354 13336 59360 13388
rect 59412 13376 59418 13388
rect 214190 13376 214196 13388
rect 59412 13348 214196 13376
rect 59412 13336 59418 13348
rect 214190 13336 214196 13348
rect 214248 13336 214254 13388
rect 243170 13336 243176 13388
rect 243228 13376 243234 13388
rect 430850 13376 430856 13388
rect 243228 13348 430856 13376
rect 243228 13336 243234 13348
rect 430850 13336 430856 13348
rect 430908 13336 430914 13388
rect 56042 13268 56048 13320
rect 56100 13308 56106 13320
rect 214374 13308 214380 13320
rect 56100 13280 214380 13308
rect 56100 13268 56106 13280
rect 214374 13268 214380 13280
rect 214432 13268 214438 13320
rect 244274 13268 244280 13320
rect 244332 13308 244338 13320
rect 440326 13308 440332 13320
rect 244332 13280 440332 13308
rect 244332 13268 244338 13280
rect 440326 13268 440332 13280
rect 440384 13268 440390 13320
rect 52546 13200 52552 13252
rect 52604 13240 52610 13252
rect 214282 13240 214288 13252
rect 52604 13212 214288 13240
rect 52604 13200 52610 13212
rect 214282 13200 214288 13212
rect 214340 13200 214346 13252
rect 244458 13200 244464 13252
rect 244516 13240 244522 13252
rect 445018 13240 445024 13252
rect 244516 13212 445024 13240
rect 244516 13200 244522 13212
rect 445018 13200 445024 13212
rect 445076 13200 445082 13252
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 210234 13172 210240 13184
rect 8812 13144 210240 13172
rect 8812 13132 8818 13144
rect 210234 13132 210240 13144
rect 210292 13132 210298 13184
rect 244366 13132 244372 13184
rect 244424 13172 244430 13184
rect 448606 13172 448612 13184
rect 244424 13144 448612 13172
rect 244424 13132 244430 13144
rect 448606 13132 448612 13144
rect 448664 13132 448670 13184
rect 3602 13064 3608 13116
rect 3660 13104 3666 13116
rect 210142 13104 210148 13116
rect 3660 13076 210148 13104
rect 3660 13064 3666 13076
rect 210142 13064 210148 13076
rect 210200 13064 210206 13116
rect 245654 13064 245660 13116
rect 245712 13104 245718 13116
rect 459186 13104 459192 13116
rect 245712 13076 459192 13104
rect 245712 13064 245718 13076
rect 459186 13064 459192 13076
rect 459244 13064 459250 13116
rect 230750 12180 230756 12232
rect 230808 12220 230814 12232
rect 264974 12220 264980 12232
rect 230808 12192 264980 12220
rect 230808 12180 230814 12192
rect 264974 12180 264980 12192
rect 265032 12180 265038 12232
rect 114738 12112 114744 12164
rect 114796 12152 114802 12164
rect 218330 12152 218336 12164
rect 114796 12124 218336 12152
rect 114796 12112 114802 12124
rect 218330 12112 218336 12124
rect 218388 12112 218394 12164
rect 236178 12112 236184 12164
rect 236236 12152 236242 12164
rect 330386 12152 330392 12164
rect 236236 12124 330392 12152
rect 236236 12112 236242 12124
rect 330386 12112 330392 12124
rect 330444 12112 330450 12164
rect 111610 12044 111616 12096
rect 111668 12084 111674 12096
rect 218238 12084 218244 12096
rect 111668 12056 218244 12084
rect 111668 12044 111674 12056
rect 218238 12044 218244 12056
rect 218296 12044 218302 12096
rect 257430 12044 257436 12096
rect 257488 12084 257494 12096
rect 415394 12084 415400 12096
rect 257488 12056 415400 12084
rect 257488 12044 257494 12056
rect 415394 12044 415400 12056
rect 415452 12044 415458 12096
rect 15930 11976 15936 12028
rect 15988 12016 15994 12028
rect 178678 12016 178684 12028
rect 15988 11988 178684 12016
rect 15988 11976 15994 11988
rect 178678 11976 178684 11988
rect 178736 11976 178742 12028
rect 178770 11976 178776 12028
rect 178828 12016 178834 12028
rect 212626 12016 212632 12028
rect 178828 11988 212632 12016
rect 178828 11976 178834 11988
rect 212626 11976 212632 11988
rect 212684 11976 212690 12028
rect 241514 11976 241520 12028
rect 241572 12016 241578 12028
rect 406010 12016 406016 12028
rect 241572 11988 406016 12016
rect 241572 11976 241578 11988
rect 406010 11976 406016 11988
rect 406068 11976 406074 12028
rect 36722 11908 36728 11960
rect 36780 11948 36786 11960
rect 212718 11948 212724 11960
rect 36780 11920 212724 11948
rect 36780 11908 36786 11920
rect 212718 11908 212724 11920
rect 212776 11908 212782 11960
rect 241606 11908 241612 11960
rect 241664 11948 241670 11960
rect 409138 11948 409144 11960
rect 241664 11920 409144 11948
rect 241664 11908 241670 11920
rect 409138 11908 409144 11920
rect 409196 11908 409202 11960
rect 33594 11840 33600 11892
rect 33652 11880 33658 11892
rect 213362 11880 213368 11892
rect 33652 11852 213368 11880
rect 33652 11840 33658 11852
rect 213362 11840 213368 11852
rect 213420 11840 213426 11892
rect 242986 11840 242992 11892
rect 243044 11880 243050 11892
rect 420178 11880 420184 11892
rect 243044 11852 420184 11880
rect 243044 11840 243050 11852
rect 420178 11840 420184 11852
rect 420236 11840 420242 11892
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 211522 11812 211528 11824
rect 26292 11784 211528 11812
rect 26292 11772 26298 11784
rect 211522 11772 211528 11784
rect 211580 11772 211586 11824
rect 243078 11772 243084 11824
rect 243136 11812 243142 11824
rect 423766 11812 423772 11824
rect 243136 11784 423772 11812
rect 243136 11772 243142 11784
rect 423766 11772 423772 11784
rect 423824 11772 423830 11824
rect 21818 11704 21824 11756
rect 21876 11744 21882 11756
rect 211246 11744 211252 11756
rect 21876 11716 211252 11744
rect 21876 11704 21882 11716
rect 211246 11704 211252 11716
rect 211304 11704 211310 11756
rect 220814 11704 220820 11756
rect 220872 11744 220878 11756
rect 221366 11744 221372 11756
rect 220872 11716 221372 11744
rect 220872 11704 220878 11716
rect 221366 11704 221372 11716
rect 221424 11704 221430 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 426802 11744 426808 11756
rect 242952 11716 426808 11744
rect 242952 11704 242958 11716
rect 426802 11704 426808 11716
rect 426860 11704 426866 11756
rect 186958 10752 186964 10804
rect 187016 10792 187022 10804
rect 218974 10792 218980 10804
rect 187016 10764 218980 10792
rect 187016 10752 187022 10764
rect 218974 10752 218980 10764
rect 219032 10752 219038 10804
rect 159358 10684 159364 10736
rect 159416 10724 159422 10736
rect 218790 10724 218796 10736
rect 159416 10696 218796 10724
rect 159416 10684 159422 10696
rect 218790 10684 218796 10696
rect 218848 10684 218854 10736
rect 97442 10616 97448 10668
rect 97500 10656 97506 10668
rect 216858 10656 216864 10668
rect 97500 10628 216864 10656
rect 97500 10616 97506 10628
rect 216858 10616 216864 10628
rect 216916 10616 216922 10668
rect 237650 10616 237656 10668
rect 237708 10656 237714 10668
rect 359458 10656 359464 10668
rect 237708 10628 359464 10656
rect 237708 10616 237714 10628
rect 359458 10616 359464 10628
rect 359516 10616 359522 10668
rect 93946 10548 93952 10600
rect 94004 10588 94010 10600
rect 217226 10588 217232 10600
rect 94004 10560 217232 10588
rect 94004 10548 94010 10560
rect 217226 10548 217232 10560
rect 217284 10548 217290 10600
rect 238846 10548 238852 10600
rect 238904 10588 238910 10600
rect 370130 10588 370136 10600
rect 238904 10560 370136 10588
rect 238904 10548 238910 10560
rect 370130 10548 370136 10560
rect 370188 10548 370194 10600
rect 89898 10480 89904 10532
rect 89956 10520 89962 10532
rect 217502 10520 217508 10532
rect 89956 10492 217508 10520
rect 89956 10480 89962 10492
rect 217502 10480 217508 10492
rect 217560 10480 217566 10532
rect 238754 10480 238760 10532
rect 238812 10520 238818 10532
rect 374086 10520 374092 10532
rect 238812 10492 374092 10520
rect 238812 10480 238818 10492
rect 374086 10480 374092 10492
rect 374144 10480 374150 10532
rect 79226 10412 79232 10464
rect 79284 10452 79290 10464
rect 215478 10452 215484 10464
rect 79284 10424 215484 10452
rect 79284 10412 79290 10424
rect 215478 10412 215484 10424
rect 215536 10412 215542 10464
rect 241422 10412 241428 10464
rect 241480 10452 241486 10464
rect 390646 10452 390652 10464
rect 241480 10424 390652 10452
rect 241480 10412 241486 10424
rect 390646 10412 390652 10424
rect 390704 10412 390710 10464
rect 75914 10344 75920 10396
rect 75972 10384 75978 10396
rect 215570 10384 215576 10396
rect 75972 10356 215576 10384
rect 75972 10344 75978 10356
rect 215570 10344 215576 10356
rect 215628 10344 215634 10396
rect 240318 10344 240324 10396
rect 240376 10384 240382 10396
rect 395338 10384 395344 10396
rect 240376 10356 395344 10384
rect 240376 10344 240382 10356
rect 395338 10344 395344 10356
rect 395396 10344 395402 10396
rect 11146 10276 11152 10328
rect 11204 10316 11210 10328
rect 188338 10316 188344 10328
rect 11204 10288 188344 10316
rect 11204 10276 11210 10288
rect 188338 10276 188344 10288
rect 188396 10276 188402 10328
rect 252738 10276 252744 10328
rect 252796 10316 252802 10328
rect 553762 10316 553768 10328
rect 252796 10288 553768 10316
rect 252796 10276 252802 10288
rect 553762 10276 553768 10288
rect 553820 10276 553826 10328
rect 125870 9392 125876 9444
rect 125928 9432 125934 9444
rect 215386 9432 215392 9444
rect 125928 9404 215392 9432
rect 125928 9392 125934 9404
rect 215386 9392 215392 9404
rect 215444 9392 215450 9444
rect 69106 9324 69112 9376
rect 69164 9364 69170 9376
rect 216214 9364 216220 9376
rect 69164 9336 216220 9364
rect 69164 9324 69170 9336
rect 216214 9324 216220 9336
rect 216272 9324 216278 9376
rect 62022 9256 62028 9308
rect 62080 9296 62086 9308
rect 214742 9296 214748 9308
rect 62080 9268 214748 9296
rect 62080 9256 62086 9268
rect 214742 9256 214748 9268
rect 214800 9256 214806 9308
rect 234798 9256 234804 9308
rect 234856 9296 234862 9308
rect 324406 9296 324412 9308
rect 234856 9268 324412 9296
rect 234856 9256 234862 9268
rect 324406 9256 324412 9268
rect 324464 9256 324470 9308
rect 58434 9188 58440 9240
rect 58492 9228 58498 9240
rect 214006 9228 214012 9240
rect 58492 9200 214012 9228
rect 58492 9188 58498 9200
rect 214006 9188 214012 9200
rect 214064 9188 214070 9240
rect 236086 9188 236092 9240
rect 236144 9228 236150 9240
rect 338666 9228 338672 9240
rect 236144 9200 338672 9228
rect 236144 9188 236150 9200
rect 338666 9188 338672 9200
rect 338724 9188 338730 9240
rect 54938 9120 54944 9172
rect 54996 9160 55002 9172
rect 214098 9160 214104 9172
rect 54996 9132 214104 9160
rect 54996 9120 55002 9132
rect 214098 9120 214104 9132
rect 214156 9120 214162 9172
rect 235994 9120 236000 9172
rect 236052 9160 236058 9172
rect 342162 9160 342168 9172
rect 236052 9132 342168 9160
rect 236052 9120 236058 9132
rect 342162 9120 342168 9132
rect 342220 9120 342226 9172
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 209958 9092 209964 9104
rect 7708 9064 209964 9092
rect 7708 9052 7714 9064
rect 209958 9052 209964 9064
rect 210016 9052 210022 9104
rect 237466 9052 237472 9104
rect 237524 9092 237530 9104
rect 349246 9092 349252 9104
rect 237524 9064 349252 9092
rect 237524 9052 237530 9064
rect 349246 9052 349252 9064
rect 349304 9052 349310 9104
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 209866 9024 209872 9036
rect 2924 8996 209872 9024
rect 2924 8984 2930 8996
rect 209866 8984 209872 8996
rect 209924 8984 209930 9036
rect 237374 8984 237380 9036
rect 237432 9024 237438 9036
rect 352834 9024 352840 9036
rect 237432 8996 352840 9024
rect 237432 8984 237438 8996
rect 352834 8984 352840 8996
rect 352892 8984 352898 9036
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 210050 8956 210056 8968
rect 1728 8928 210056 8956
rect 1728 8916 1734 8928
rect 210050 8916 210056 8928
rect 210108 8916 210114 8968
rect 237558 8916 237564 8968
rect 237616 8956 237622 8968
rect 356330 8956 356336 8968
rect 237616 8928 356336 8956
rect 237616 8916 237622 8928
rect 356330 8916 356336 8928
rect 356388 8916 356394 8968
rect 158898 7896 158904 7948
rect 158956 7936 158962 7948
rect 222654 7936 222660 7948
rect 158956 7908 222660 7936
rect 158956 7896 158962 7908
rect 222654 7896 222660 7908
rect 222712 7896 222718 7948
rect 233326 7896 233332 7948
rect 233384 7936 233390 7948
rect 303154 7936 303160 7948
rect 233384 7908 303160 7936
rect 233384 7896 233390 7908
rect 303154 7896 303160 7908
rect 303212 7896 303218 7948
rect 155402 7828 155408 7880
rect 155460 7868 155466 7880
rect 220078 7868 220084 7880
rect 155460 7840 220084 7868
rect 155460 7828 155466 7840
rect 220078 7828 220084 7840
rect 220136 7828 220142 7880
rect 233234 7828 233240 7880
rect 233292 7868 233298 7880
rect 306742 7868 306748 7880
rect 233292 7840 306748 7868
rect 233292 7828 233298 7840
rect 306742 7828 306748 7840
rect 306800 7828 306806 7880
rect 151906 7760 151912 7812
rect 151964 7800 151970 7812
rect 220998 7800 221004 7812
rect 151964 7772 221004 7800
rect 151964 7760 151970 7772
rect 220998 7760 221004 7772
rect 221056 7760 221062 7812
rect 234614 7760 234620 7812
rect 234672 7800 234678 7812
rect 317322 7800 317328 7812
rect 234672 7772 317328 7800
rect 234672 7760 234678 7772
rect 317322 7760 317328 7772
rect 317380 7760 317386 7812
rect 148318 7692 148324 7744
rect 148376 7732 148382 7744
rect 221182 7732 221188 7744
rect 148376 7704 221188 7732
rect 148376 7692 148382 7704
rect 221182 7692 221188 7704
rect 221240 7692 221246 7744
rect 235902 7692 235908 7744
rect 235960 7732 235966 7744
rect 320910 7732 320916 7744
rect 235960 7704 320916 7732
rect 235960 7692 235966 7704
rect 320910 7692 320916 7704
rect 320968 7692 320974 7744
rect 144730 7624 144736 7676
rect 144788 7664 144794 7676
rect 221090 7664 221096 7676
rect 144788 7636 221096 7664
rect 144788 7624 144794 7636
rect 221090 7624 221096 7636
rect 221148 7624 221154 7676
rect 248506 7624 248512 7676
rect 248564 7664 248570 7676
rect 492306 7664 492312 7676
rect 248564 7636 492312 7664
rect 248564 7624 248570 7636
rect 492306 7624 492312 7636
rect 492364 7624 492370 7676
rect 141234 7556 141240 7608
rect 141292 7596 141298 7608
rect 221274 7596 221280 7608
rect 141292 7568 221280 7596
rect 141292 7556 141298 7568
rect 221274 7556 221280 7568
rect 221332 7556 221338 7608
rect 251450 7556 251456 7608
rect 251508 7596 251514 7608
rect 529014 7596 529020 7608
rect 251508 7568 529020 7596
rect 251508 7556 251514 7568
rect 529014 7556 529020 7568
rect 529072 7556 529078 7608
rect 197906 6468 197912 6520
rect 197964 6508 197970 6520
rect 225138 6508 225144 6520
rect 197964 6480 225144 6508
rect 197964 6468 197970 6480
rect 225138 6468 225144 6480
rect 225196 6468 225202 6520
rect 231854 6468 231860 6520
rect 231912 6508 231918 6520
rect 285398 6508 285404 6520
rect 231912 6480 285404 6508
rect 231912 6468 231918 6480
rect 285398 6468 285404 6480
rect 285456 6468 285462 6520
rect 187326 6400 187332 6452
rect 187384 6440 187390 6452
rect 223942 6440 223948 6452
rect 187384 6412 223948 6440
rect 187384 6400 187390 6412
rect 223942 6400 223948 6412
rect 224000 6400 224006 6452
rect 240134 6400 240140 6452
rect 240192 6440 240198 6452
rect 388254 6440 388260 6452
rect 240192 6412 388260 6440
rect 240192 6400 240198 6412
rect 388254 6400 388260 6412
rect 388312 6400 388318 6452
rect 183738 6332 183744 6384
rect 183796 6372 183802 6384
rect 223850 6372 223856 6384
rect 183796 6344 223856 6372
rect 183796 6332 183802 6344
rect 223850 6332 223856 6344
rect 223908 6332 223914 6384
rect 256326 6332 256332 6384
rect 256384 6372 256390 6384
rect 562042 6372 562048 6384
rect 256384 6344 562048 6372
rect 256384 6332 256390 6344
rect 562042 6332 562048 6344
rect 562100 6332 562106 6384
rect 180242 6264 180248 6316
rect 180300 6304 180306 6316
rect 223758 6304 223764 6316
rect 180300 6276 223764 6304
rect 180300 6264 180306 6276
rect 223758 6264 223764 6276
rect 223816 6264 223822 6316
rect 254026 6264 254032 6316
rect 254084 6304 254090 6316
rect 566826 6304 566832 6316
rect 254084 6276 566832 6304
rect 254084 6264 254090 6276
rect 566826 6264 566832 6276
rect 566884 6264 566890 6316
rect 128170 6196 128176 6248
rect 128228 6236 128234 6248
rect 219802 6236 219808 6248
rect 128228 6208 219808 6236
rect 128228 6196 128234 6208
rect 219802 6196 219808 6208
rect 219860 6196 219866 6248
rect 253934 6196 253940 6248
rect 253992 6236 253998 6248
rect 569126 6236 569132 6248
rect 253992 6208 569132 6236
rect 253992 6196 253998 6208
rect 569126 6196 569132 6208
rect 569184 6196 569190 6248
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 209038 6168 209044 6180
rect 6512 6140 209044 6168
rect 6512 6128 6518 6140
rect 209038 6128 209044 6140
rect 209096 6128 209102 6180
rect 254118 6128 254124 6180
rect 254176 6168 254182 6180
rect 572714 6168 572720 6180
rect 254176 6140 572720 6168
rect 254176 6128 254182 6140
rect 572714 6128 572720 6140
rect 572772 6128 572778 6180
rect 201586 5380 201592 5432
rect 201644 5420 201650 5432
rect 225506 5420 225512 5432
rect 201644 5392 225512 5420
rect 201644 5380 201650 5392
rect 225506 5380 225512 5392
rect 225564 5380 225570 5432
rect 176746 5312 176752 5364
rect 176804 5352 176810 5364
rect 224402 5352 224408 5364
rect 176804 5324 224408 5352
rect 176804 5312 176810 5324
rect 224402 5312 224408 5324
rect 224460 5312 224466 5364
rect 169570 5244 169576 5296
rect 169628 5284 169634 5296
rect 222562 5284 222568 5296
rect 169628 5256 222568 5284
rect 169628 5244 169634 5256
rect 222562 5244 222568 5256
rect 222620 5244 222626 5296
rect 166074 5176 166080 5228
rect 166132 5216 166138 5228
rect 223482 5216 223488 5228
rect 166132 5188 223488 5216
rect 166132 5176 166138 5188
rect 223482 5176 223488 5188
rect 223540 5176 223546 5228
rect 230658 5176 230664 5228
rect 230716 5216 230722 5228
rect 262950 5216 262956 5228
rect 230716 5188 262956 5216
rect 230716 5176 230722 5188
rect 262950 5176 262956 5188
rect 263008 5176 263014 5228
rect 162486 5108 162492 5160
rect 162544 5148 162550 5160
rect 222378 5148 222384 5160
rect 162544 5120 222384 5148
rect 162544 5108 162550 5120
rect 222378 5108 222384 5120
rect 222436 5108 222442 5160
rect 249794 5108 249800 5160
rect 249852 5148 249858 5160
rect 519538 5148 519544 5160
rect 249852 5120 519544 5148
rect 249852 5108 249858 5120
rect 519538 5108 519544 5120
rect 519596 5108 519602 5160
rect 157794 5040 157800 5092
rect 157852 5080 157858 5092
rect 222470 5080 222476 5092
rect 157852 5052 222476 5080
rect 157852 5040 157858 5052
rect 222470 5040 222476 5052
rect 222528 5040 222534 5092
rect 251358 5040 251364 5092
rect 251416 5080 251422 5092
rect 525426 5080 525432 5092
rect 251416 5052 525432 5080
rect 251416 5040 251422 5052
rect 525426 5040 525432 5052
rect 525484 5040 525490 5092
rect 150618 4972 150624 5024
rect 150676 5012 150682 5024
rect 220906 5012 220912 5024
rect 150676 4984 220912 5012
rect 150676 4972 150682 4984
rect 220906 4972 220912 4984
rect 220964 4972 220970 5024
rect 251266 4972 251272 5024
rect 251324 5012 251330 5024
rect 533706 5012 533712 5024
rect 251324 4984 533712 5012
rect 251324 4972 251330 4984
rect 533706 4972 533712 4984
rect 533764 4972 533770 5024
rect 143534 4904 143540 4956
rect 143592 4944 143598 4956
rect 221642 4944 221648 4956
rect 143592 4916 221648 4944
rect 143592 4904 143598 4916
rect 221642 4904 221648 4916
rect 221700 4904 221706 4956
rect 251174 4904 251180 4956
rect 251232 4944 251238 4956
rect 537202 4944 537208 4956
rect 251232 4916 537208 4944
rect 251232 4904 251238 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 126974 4836 126980 4888
rect 127032 4876 127038 4888
rect 219710 4876 219716 4888
rect 127032 4848 219716 4876
rect 127032 4836 127038 4848
rect 219710 4836 219716 4848
rect 219768 4836 219774 4888
rect 229370 4836 229376 4888
rect 229428 4876 229434 4888
rect 247586 4876 247592 4888
rect 229428 4848 247592 4876
rect 229428 4836 229434 4848
rect 247586 4836 247592 4848
rect 247644 4836 247650 4888
rect 252646 4836 252652 4888
rect 252704 4876 252710 4888
rect 547874 4876 547880 4888
rect 252704 4848 547880 4876
rect 252704 4836 252710 4848
rect 547874 4836 547880 4848
rect 547932 4836 547938 4888
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 203518 4808 203524 4820
rect 19484 4780 203524 4808
rect 19484 4768 19490 4780
rect 203518 4768 203524 4780
rect 203576 4768 203582 4820
rect 205082 4768 205088 4820
rect 205140 4808 205146 4820
rect 225782 4808 225788 4820
rect 205140 4780 225788 4808
rect 205140 4768 205146 4780
rect 225782 4768 225788 4780
rect 225840 4768 225846 4820
rect 229462 4768 229468 4820
rect 229520 4808 229526 4820
rect 252370 4808 252376 4820
rect 229520 4780 252376 4808
rect 229520 4768 229526 4780
rect 252370 4768 252376 4780
rect 252428 4768 252434 4820
rect 252554 4768 252560 4820
rect 252612 4808 252618 4820
rect 554958 4808 554964 4820
rect 252612 4780 554964 4808
rect 252612 4768 252618 4780
rect 554958 4768 554964 4780
rect 555016 4768 555022 4820
rect 230566 4156 230572 4208
rect 230624 4196 230630 4208
rect 230624 4168 234660 4196
rect 230624 4156 230630 4168
rect 186130 4088 186136 4140
rect 186188 4128 186194 4140
rect 224310 4128 224316 4140
rect 186188 4100 224316 4128
rect 186188 4088 186194 4100
rect 224310 4088 224316 4100
rect 224368 4088 224374 4140
rect 227898 4088 227904 4140
rect 227956 4128 227962 4140
rect 229830 4128 229836 4140
rect 227956 4100 229836 4128
rect 227956 4088 227962 4100
rect 229830 4088 229836 4100
rect 229888 4088 229894 4140
rect 234632 4128 234660 4168
rect 234632 4100 238754 4128
rect 182542 4020 182548 4072
rect 182600 4060 182606 4072
rect 209130 4060 209136 4072
rect 182600 4032 209136 4060
rect 182600 4020 182606 4032
rect 209130 4020 209136 4032
rect 209188 4020 209194 4072
rect 210970 4020 210976 4072
rect 211028 4060 211034 4072
rect 227162 4060 227168 4072
rect 211028 4032 227168 4060
rect 211028 4020 211034 4032
rect 227162 4020 227168 4032
rect 227220 4020 227226 4072
rect 95142 3952 95148 4004
rect 95200 3992 95206 4004
rect 141418 3992 141424 4004
rect 95200 3964 141424 3992
rect 95200 3952 95206 3964
rect 141418 3952 141424 3964
rect 141476 3952 141482 4004
rect 151814 3952 151820 4004
rect 151872 3992 151878 4004
rect 153010 3992 153016 4004
rect 151872 3964 153016 3992
rect 151872 3952 151878 3964
rect 153010 3952 153016 3964
rect 153068 3952 153074 4004
rect 168374 3952 168380 4004
rect 168432 3992 168438 4004
rect 207658 3992 207664 4004
rect 168432 3964 207664 3992
rect 168432 3952 168438 3964
rect 207658 3952 207664 3964
rect 207716 3952 207722 4004
rect 213362 3952 213368 4004
rect 213420 3992 213426 4004
rect 226518 3992 226524 4004
rect 213420 3964 226524 3992
rect 213420 3952 213426 3964
rect 226518 3952 226524 3964
rect 226576 3952 226582 4004
rect 104526 3884 104532 3936
rect 104584 3924 104590 3936
rect 159358 3924 159364 3936
rect 104584 3896 159364 3924
rect 104584 3884 104590 3896
rect 159358 3884 159364 3896
rect 159416 3884 159422 3936
rect 164878 3884 164884 3936
rect 164936 3924 164942 3936
rect 213178 3924 213184 3936
rect 164936 3896 213184 3924
rect 164936 3884 164942 3896
rect 213178 3884 213184 3896
rect 213236 3884 213242 3936
rect 215662 3884 215668 3936
rect 215720 3924 215726 3936
rect 225598 3924 225604 3936
rect 215720 3896 225604 3924
rect 215720 3884 215726 3896
rect 225598 3884 225604 3896
rect 225656 3884 225662 3936
rect 99834 3816 99840 3868
rect 99892 3856 99898 3868
rect 155218 3856 155224 3868
rect 99892 3828 155224 3856
rect 99892 3816 99898 3828
rect 155218 3816 155224 3828
rect 155276 3816 155282 3868
rect 167178 3816 167184 3868
rect 167236 3856 167242 3868
rect 215938 3856 215944 3868
rect 167236 3828 215944 3856
rect 167236 3816 167242 3828
rect 215938 3816 215944 3828
rect 215996 3816 216002 3868
rect 219250 3816 219256 3868
rect 219308 3856 219314 3868
rect 222838 3856 222844 3868
rect 219308 3828 222844 3856
rect 219308 3816 219314 3828
rect 222838 3816 222844 3828
rect 222896 3816 222902 3868
rect 238726 3856 238754 4100
rect 256234 4088 256240 4140
rect 256292 4128 256298 4140
rect 259454 4128 259460 4140
rect 256292 4100 259460 4128
rect 256292 4088 256298 4100
rect 259454 4088 259460 4100
rect 259512 4088 259518 4140
rect 261754 3856 261760 3868
rect 238726 3828 261760 3856
rect 261754 3816 261760 3828
rect 261812 3816 261818 3868
rect 276014 3816 276020 3868
rect 276072 3856 276078 3868
rect 276750 3856 276756 3868
rect 276072 3828 276756 3856
rect 276072 3816 276078 3828
rect 276750 3816 276756 3828
rect 276808 3816 276814 3868
rect 299566 3816 299572 3868
rect 299624 3856 299630 3868
rect 300762 3856 300768 3868
rect 299624 3828 300768 3856
rect 299624 3816 299630 3828
rect 300762 3816 300768 3828
rect 300820 3816 300826 3868
rect 418798 3816 418804 3868
rect 418856 3856 418862 3868
rect 580994 3856 581000 3868
rect 418856 3828 581000 3856
rect 418856 3816 418862 3828
rect 580994 3816 581000 3828
rect 581052 3816 581058 3868
rect 77386 3748 77392 3800
rect 77444 3788 77450 3800
rect 133138 3788 133144 3800
rect 77444 3760 133144 3788
rect 77444 3748 77450 3760
rect 133138 3748 133144 3760
rect 133196 3748 133202 3800
rect 136450 3748 136456 3800
rect 136508 3788 136514 3800
rect 213270 3788 213276 3800
rect 136508 3760 213276 3788
rect 136508 3748 136514 3760
rect 213270 3748 213276 3760
rect 213328 3748 213334 3800
rect 214466 3748 214472 3800
rect 214524 3788 214530 3800
rect 226886 3788 226892 3800
rect 214524 3760 226892 3788
rect 214524 3748 214530 3760
rect 226886 3748 226892 3760
rect 226944 3748 226950 3800
rect 256050 3748 256056 3800
rect 256108 3788 256114 3800
rect 465166 3788 465172 3800
rect 256108 3760 465172 3788
rect 256108 3748 256114 3760
rect 465166 3748 465172 3760
rect 465224 3748 465230 3800
rect 470566 3760 480254 3788
rect 108114 3680 108120 3732
rect 108172 3720 108178 3732
rect 186958 3720 186964 3732
rect 108172 3692 186964 3720
rect 108172 3680 108178 3692
rect 186958 3680 186964 3692
rect 187016 3680 187022 3732
rect 196802 3680 196808 3732
rect 196860 3720 196866 3732
rect 210418 3720 210424 3732
rect 196860 3692 210424 3720
rect 196860 3680 196866 3692
rect 210418 3680 210424 3692
rect 210476 3680 210482 3732
rect 212166 3680 212172 3732
rect 212224 3720 212230 3732
rect 226610 3720 226616 3732
rect 212224 3692 226616 3720
rect 212224 3680 212230 3692
rect 226610 3680 226616 3692
rect 226668 3680 226674 3732
rect 228082 3680 228088 3732
rect 228140 3720 228146 3732
rect 235810 3720 235816 3732
rect 228140 3692 235816 3720
rect 228140 3680 228146 3692
rect 235810 3680 235816 3692
rect 235868 3680 235874 3732
rect 257338 3680 257344 3732
rect 257396 3720 257402 3732
rect 468662 3720 468668 3732
rect 257396 3692 468668 3720
rect 257396 3680 257402 3692
rect 468662 3680 468668 3692
rect 468720 3680 468726 3732
rect 132954 3612 132960 3664
rect 133012 3652 133018 3664
rect 219618 3652 219624 3664
rect 133012 3624 219624 3652
rect 133012 3612 133018 3624
rect 219618 3612 219624 3624
rect 219676 3612 219682 3664
rect 227806 3612 227812 3664
rect 227864 3652 227870 3664
rect 237006 3652 237012 3664
rect 227864 3624 237012 3652
rect 227864 3612 227870 3624
rect 237006 3612 237012 3624
rect 237064 3612 237070 3664
rect 237374 3612 237380 3664
rect 237432 3652 237438 3664
rect 258258 3652 258264 3664
rect 237432 3624 258264 3652
rect 237432 3612 237438 3624
rect 258258 3612 258264 3624
rect 258316 3612 258322 3664
rect 258718 3612 258724 3664
rect 258776 3652 258782 3664
rect 470566 3652 470594 3760
rect 479334 3720 479340 3732
rect 258776 3624 470594 3652
rect 473188 3692 479340 3720
rect 258776 3612 258782 3624
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 125870 3584 125876 3596
rect 72660 3556 125876 3584
rect 72660 3544 72666 3556
rect 125870 3544 125876 3556
rect 125928 3544 125934 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 219526 3584 219532 3596
rect 129424 3556 219532 3584
rect 129424 3544 129430 3556
rect 219526 3544 219532 3556
rect 219584 3544 219590 3596
rect 230106 3544 230112 3596
rect 230164 3584 230170 3596
rect 244090 3584 244096 3596
rect 230164 3556 244096 3584
rect 230164 3544 230170 3556
rect 244090 3544 244096 3556
rect 244148 3544 244154 3596
rect 248414 3544 248420 3596
rect 248472 3584 248478 3596
rect 248472 3556 253612 3584
rect 248472 3544 248478 3556
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 44266 3476 44272 3528
rect 44324 3516 44330 3528
rect 44324 3488 175044 3516
rect 44324 3476 44330 3488
rect 52454 3408 52460 3460
rect 52512 3448 52518 3460
rect 53374 3448 53380 3460
rect 52512 3420 53380 3448
rect 52512 3408 52518 3420
rect 53374 3408 53380 3420
rect 53432 3408 53438 3460
rect 175016 3448 175044 3488
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177850 3516 177856 3528
rect 176712 3488 177856 3516
rect 176712 3476 176718 3488
rect 177850 3476 177856 3488
rect 177908 3476 177914 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202690 3516 202696 3528
rect 201552 3488 202696 3516
rect 201552 3476 201558 3488
rect 202690 3476 202696 3488
rect 202748 3476 202754 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 226426 3516 226432 3528
rect 224000 3488 226432 3516
rect 224000 3476 224006 3488
rect 226426 3476 226432 3488
rect 226484 3476 226490 3528
rect 227530 3476 227536 3528
rect 227588 3516 227594 3528
rect 227990 3516 227996 3528
rect 227588 3488 227996 3516
rect 227588 3476 227594 3488
rect 227990 3476 227996 3488
rect 228048 3476 228054 3528
rect 231118 3476 231124 3528
rect 231176 3516 231182 3528
rect 232222 3516 232228 3528
rect 231176 3488 232228 3516
rect 231176 3476 231182 3488
rect 232222 3476 232228 3488
rect 232280 3476 232286 3528
rect 232332 3488 238754 3516
rect 178770 3448 178776 3460
rect 55186 3420 161474 3448
rect 175016 3420 178776 3448
rect 47854 3340 47860 3392
rect 47912 3380 47918 3392
rect 55186 3380 55214 3420
rect 47912 3352 55214 3380
rect 47912 3340 47918 3352
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 20622 3272 20628 3324
rect 20680 3312 20686 3324
rect 25498 3312 25504 3324
rect 20680 3284 25504 3312
rect 20680 3272 20686 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 161446 3312 161474 3420
rect 178770 3408 178776 3420
rect 178828 3408 178834 3460
rect 207750 3448 207756 3460
rect 180766 3420 207756 3448
rect 180766 3312 180794 3420
rect 207750 3408 207756 3420
rect 207808 3408 207814 3460
rect 229186 3408 229192 3460
rect 229244 3448 229250 3460
rect 232332 3448 232360 3488
rect 229244 3420 232360 3448
rect 238726 3448 238754 3488
rect 250438 3476 250444 3528
rect 250496 3516 250502 3528
rect 251174 3516 251180 3528
rect 250496 3488 251180 3516
rect 250496 3476 250502 3488
rect 251174 3476 251180 3488
rect 251232 3476 251238 3528
rect 253474 3448 253480 3460
rect 238726 3420 253480 3448
rect 229244 3408 229250 3420
rect 253474 3408 253480 3420
rect 253532 3408 253538 3460
rect 253584 3448 253612 3556
rect 256142 3544 256148 3596
rect 256200 3584 256206 3596
rect 473188 3584 473216 3692
rect 479334 3680 479340 3692
rect 479392 3680 479398 3732
rect 480226 3652 480254 3760
rect 480530 3652 480536 3664
rect 480226 3624 480536 3652
rect 480530 3612 480536 3624
rect 480588 3612 480594 3664
rect 256200 3556 473216 3584
rect 256200 3544 256206 3556
rect 473354 3544 473360 3596
rect 473412 3584 473418 3596
rect 474182 3584 474188 3596
rect 473412 3556 474188 3584
rect 473412 3544 473418 3556
rect 474182 3544 474188 3556
rect 474240 3544 474246 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482462 3584 482468 3596
rect 481692 3556 482468 3584
rect 481692 3544 481698 3556
rect 482462 3544 482468 3556
rect 482520 3544 482526 3596
rect 255958 3476 255964 3528
rect 256016 3516 256022 3528
rect 491110 3516 491116 3528
rect 256016 3488 491116 3516
rect 256016 3476 256022 3488
rect 491110 3476 491116 3488
rect 491168 3476 491174 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 501782 3448 501788 3460
rect 253584 3420 501788 3448
rect 501782 3408 501788 3420
rect 501840 3408 501846 3460
rect 229278 3340 229284 3392
rect 229336 3380 229342 3392
rect 246390 3380 246396 3392
rect 229336 3352 246396 3380
rect 229336 3340 229342 3352
rect 246390 3340 246396 3352
rect 246448 3340 246454 3392
rect 249978 3340 249984 3392
rect 250036 3380 250042 3392
rect 256694 3380 256700 3392
rect 250036 3352 256700 3380
rect 250036 3340 250042 3352
rect 256694 3340 256700 3352
rect 256752 3340 256758 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365806 3340 365812 3392
rect 365864 3380 365870 3392
rect 367002 3380 367008 3392
rect 365864 3352 367008 3380
rect 365864 3340 365870 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 161446 3284 180794 3312
rect 226334 3136 226340 3188
rect 226392 3176 226398 3188
rect 228174 3176 228180 3188
rect 226392 3148 228180 3176
rect 226392 3136 226398 3148
rect 228174 3136 228180 3148
rect 228232 3136 228238 3188
rect 242158 3136 242164 3188
rect 242216 3176 242222 3188
rect 245194 3176 245200 3188
rect 242216 3148 245200 3176
rect 242216 3136 242222 3148
rect 245194 3136 245200 3148
rect 245252 3136 245258 3188
rect 232498 3068 232504 3120
rect 232556 3108 232562 3120
rect 238110 3108 238116 3120
rect 232556 3080 238116 3108
rect 232556 3068 232562 3080
rect 238110 3068 238116 3080
rect 238168 3068 238174 3120
rect 423674 960 423680 1012
rect 423732 1000 423738 1012
rect 424962 1000 424968 1012
rect 423732 972 424968 1000
rect 423732 960 423738 972
rect 424962 960 424968 972
rect 425020 960 425026 1012
rect 448514 960 448520 1012
rect 448572 1000 448578 1012
rect 449802 1000 449808 1012
rect 448572 972 449808 1000
rect 448572 960 448578 972
rect 449802 960 449808 972
rect 449860 960 449866 1012
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 405004 700544 405056 700596
rect 413652 700544 413704 700596
rect 154120 700476 154172 700528
rect 182824 700476 182876 700528
rect 296076 700476 296128 700528
rect 300124 700476 300176 700528
rect 409144 700476 409196 700528
rect 429844 700476 429896 700528
rect 137836 700408 137888 700460
rect 178684 700408 178736 700460
rect 188896 700408 188948 700460
rect 202788 700408 202840 700460
rect 293224 700408 293276 700460
rect 332508 700408 332560 700460
rect 403624 700408 403676 700460
rect 462320 700408 462372 700460
rect 105452 700340 105504 700392
rect 174544 700340 174596 700392
rect 188988 700340 189040 700392
rect 218980 700340 219032 700392
rect 291844 700340 291896 700392
rect 348792 700340 348844 700392
rect 399484 700340 399536 700392
rect 478512 700340 478564 700392
rect 89168 700272 89220 700324
rect 184204 700272 184256 700324
rect 188804 700272 188856 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 281540 700272 281592 700324
rect 295984 700272 296036 700324
rect 364984 700272 365036 700324
rect 406384 700272 406436 700324
rect 494796 700272 494848 700324
rect 509884 700272 509936 700324
rect 559656 700272 559708 700324
rect 170312 699660 170364 699712
rect 171784 699660 171836 699712
rect 395344 699660 395396 699712
rect 397460 699660 397512 699712
rect 286324 696940 286376 696992
rect 580172 696940 580224 696992
rect 508504 670692 508556 670744
rect 580172 670692 580224 670744
rect 512644 643084 512696 643136
rect 580172 643084 580224 643136
rect 501604 630640 501656 630692
rect 579988 630640 580040 630692
rect 504364 616836 504416 616888
rect 580172 616836 580224 616888
rect 297364 600244 297416 600296
rect 297824 600244 297876 600296
rect 78128 599972 78180 600024
rect 187240 599972 187292 600024
rect 297824 599972 297876 600024
rect 408040 599972 408092 600024
rect 78036 599904 78088 599956
rect 187148 599904 187200 599956
rect 78588 599836 78640 599888
rect 187332 599836 187384 599888
rect 78220 599768 78272 599820
rect 186872 599768 186924 599820
rect 78404 599700 78456 599752
rect 187056 599700 187108 599752
rect 78496 599632 78548 599684
rect 186964 599632 187016 599684
rect 297916 598884 297968 598936
rect 407948 598884 408000 598936
rect 297456 598816 297508 598868
rect 408132 598816 408184 598868
rect 297548 598748 297600 598800
rect 407580 598748 407632 598800
rect 297272 598000 297324 598052
rect 297916 598000 297968 598052
rect 102876 597252 102928 597304
rect 212448 597252 212500 597304
rect 284300 597252 284352 597304
rect 325792 597252 325844 597304
rect 434720 597252 434772 597304
rect 106096 597184 106148 597236
rect 215944 597184 215996 597236
rect 319444 597184 319496 597236
rect 427820 597184 427872 597236
rect 103428 597116 103480 597168
rect 213828 597116 213880 597168
rect 318340 597116 318392 597168
rect 426440 597116 426492 597168
rect 104808 597048 104860 597100
rect 214840 597048 214892 597100
rect 319260 597048 319312 597100
rect 320088 597048 320140 597100
rect 429200 597048 429252 597100
rect 100668 596980 100720 597032
rect 210056 596980 210108 597032
rect 211068 596980 211120 597032
rect 320916 596980 320968 597032
rect 430580 596980 430632 597032
rect 97908 596912 97960 596964
rect 207112 596912 207164 596964
rect 324412 596912 324464 596964
rect 434720 596912 434772 596964
rect 99288 596844 99340 596896
rect 208400 596844 208452 596896
rect 212448 596844 212500 596896
rect 284576 596844 284628 596896
rect 321560 596844 321612 596896
rect 322296 596844 322348 596896
rect 431960 596844 432012 596896
rect 102048 596776 102100 596828
rect 140688 596504 140740 596556
rect 172244 596504 172296 596556
rect 214840 596776 214892 596828
rect 284392 596776 284444 596828
rect 299204 596776 299256 596828
rect 313280 596776 313332 596828
rect 322940 596776 322992 596828
rect 433340 596776 433392 596828
rect 280988 596708 281040 596760
rect 318340 596708 318392 596760
rect 215944 596640 215996 596692
rect 284300 596640 284352 596692
rect 299296 596640 299348 596692
rect 314660 596640 314712 596692
rect 283104 596572 283156 596624
rect 319260 596572 319312 596624
rect 211160 596504 211212 596556
rect 283012 596504 283064 596556
rect 320916 596504 320968 596556
rect 408132 596504 408184 596556
rect 422576 596504 422628 596556
rect 136548 596436 136600 596488
rect 173348 596436 173400 596488
rect 213828 596436 213880 596488
rect 284484 596436 284536 596488
rect 284576 596436 284628 596488
rect 321560 596436 321612 596488
rect 408040 596436 408092 596488
rect 423680 596436 423732 596488
rect 131028 596368 131080 596420
rect 171876 596368 171928 596420
rect 208400 596368 208452 596420
rect 281632 596368 281684 596420
rect 319444 596368 319496 596420
rect 407948 596368 408000 596420
rect 425060 596368 425112 596420
rect 79876 596300 79928 596352
rect 92480 596300 92532 596352
rect 126888 596300 126940 596352
rect 173164 596300 173216 596352
rect 188620 596300 188672 596352
rect 202880 596300 202932 596352
rect 211068 596300 211120 596352
rect 283104 596300 283156 596352
rect 284484 596300 284536 596352
rect 322940 596300 322992 596352
rect 406476 596300 406528 596352
rect 434720 596300 434772 596352
rect 79784 596232 79836 596284
rect 94044 596232 94096 596284
rect 121368 596232 121420 596284
rect 171968 596232 172020 596284
rect 188712 596232 188764 596284
rect 204352 596232 204404 596284
rect 284392 596232 284444 596284
rect 324412 596232 324464 596284
rect 409328 596232 409380 596284
rect 444380 596232 444432 596284
rect 79968 596164 80020 596216
rect 95240 596164 95292 596216
rect 115848 596164 115900 596216
rect 172152 596164 172204 596216
rect 188528 596164 188580 596216
rect 204260 596164 204312 596216
rect 207112 596164 207164 596216
rect 280988 596164 281040 596216
rect 299388 596164 299440 596216
rect 311900 596164 311952 596216
rect 409236 596164 409288 596216
rect 455420 596164 455472 596216
rect 282184 592628 282236 592680
rect 440240 592628 440292 592680
rect 284944 590656 284996 590708
rect 580172 590656 580224 590708
rect 289084 589908 289136 589960
rect 329840 589908 329892 589960
rect 287704 588616 287756 588668
rect 324320 588616 324372 588668
rect 282276 588548 282328 588600
rect 449900 588548 449952 588600
rect 78312 587120 78364 587172
rect 186780 587120 186832 587172
rect 286416 587120 286468 587172
rect 360200 587120 360252 587172
rect 298836 585828 298888 585880
rect 354680 585828 354732 585880
rect 298008 585760 298060 585812
rect 407672 585760 407724 585812
rect 297180 585148 297232 585200
rect 298008 585148 298060 585200
rect 293316 584400 293368 584452
rect 349160 584400 349212 584452
rect 283564 582972 283616 583024
rect 339500 582972 339552 583024
rect 226248 581612 226300 581664
rect 281724 581612 281776 581664
rect 289176 581612 289228 581664
rect 345020 581612 345072 581664
rect 251088 580524 251140 580576
rect 282092 580524 282144 580576
rect 245568 580456 245620 580508
rect 281080 580456 281132 580508
rect 241428 580388 241480 580440
rect 281816 580388 281868 580440
rect 190000 580320 190052 580372
rect 215300 580320 215352 580372
rect 235908 580320 235960 580372
rect 281908 580320 281960 580372
rect 285036 580320 285088 580372
rect 335360 580320 335412 580372
rect 106188 580252 106240 580304
rect 172060 580252 172112 580304
rect 189908 580252 189960 580304
rect 219440 580252 219492 580304
rect 231768 580252 231820 580304
rect 282000 580252 282052 580304
rect 282368 580252 282420 580304
rect 459560 580252 459612 580304
rect 516784 576852 516836 576904
rect 580172 576852 580224 576904
rect 3332 565836 3384 565888
rect 32404 565836 32456 565888
rect 507124 563048 507176 563100
rect 580172 563048 580224 563100
rect 3148 553392 3200 553444
rect 22744 553392 22796 553444
rect 511264 536800 511316 536852
rect 579896 536800 579948 536852
rect 3332 527144 3384 527196
rect 14464 527144 14516 527196
rect 293868 527008 293920 527060
rect 297272 527008 297324 527060
rect 298008 527008 298060 527060
rect 187332 525784 187384 525836
rect 187700 525784 187752 525836
rect 514024 524424 514076 524476
rect 580172 524424 580224 524476
rect 502984 510620 503036 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 10324 500964 10376 501016
rect 287796 498788 287848 498840
rect 297088 498788 297140 498840
rect 78496 489812 78548 489864
rect 187700 489812 187752 489864
rect 78312 489744 78364 489796
rect 187516 489744 187568 489796
rect 297640 489744 297692 489796
rect 407764 489812 407816 489864
rect 78128 489676 78180 489728
rect 187148 489676 187200 489728
rect 77760 489608 77812 489660
rect 187332 489608 187384 489660
rect 78036 489540 78088 489592
rect 187056 489540 187108 489592
rect 78404 489472 78456 489524
rect 186964 489472 187016 489524
rect 77852 489404 77904 489456
rect 186872 489404 186924 489456
rect 78588 489336 78640 489388
rect 186780 489336 186832 489388
rect 173348 489200 173400 489252
rect 253572 489200 253624 489252
rect 218060 489132 218112 489184
rect 405004 489132 405056 489184
rect 186872 488656 186924 488708
rect 187608 488656 187660 488708
rect 187056 488588 187108 488640
rect 187424 488588 187476 488640
rect 186964 488520 187016 488572
rect 187240 488520 187292 488572
rect 79876 488452 79928 488504
rect 92940 488452 92992 488504
rect 188620 488452 188672 488504
rect 407948 488452 408000 488504
rect 425060 488452 425112 488504
rect 79784 488384 79836 488436
rect 94228 488384 94280 488436
rect 188528 488384 188580 488436
rect 204444 488384 204496 488436
rect 291936 488384 291988 488436
rect 297824 488384 297876 488436
rect 407856 488384 407908 488436
rect 408040 488384 408092 488436
rect 423680 488384 423732 488436
rect 79968 488316 80020 488368
rect 95332 488316 95384 488368
rect 297272 488316 297324 488368
rect 407488 488316 407540 488368
rect 408132 488316 408184 488368
rect 422576 488316 422628 488368
rect 299204 488248 299256 488300
rect 314292 488248 314344 488300
rect 408040 488248 408092 488300
rect 188620 488180 188672 488232
rect 202880 488180 202932 488232
rect 299296 488180 299348 488232
rect 315396 488180 315448 488232
rect 407948 488180 408000 488232
rect 188712 488112 188764 488164
rect 204904 488112 204956 488164
rect 297916 488112 297968 488164
rect 408316 488112 408368 488164
rect 188804 488044 188856 488096
rect 220084 488044 220136 488096
rect 104808 487976 104860 488028
rect 214840 487976 214892 488028
rect 230572 487976 230624 488028
rect 287796 487976 287848 488028
rect 103428 487908 103480 487960
rect 213736 487908 213788 487960
rect 219808 487908 219860 487960
rect 281540 487908 281592 487960
rect 105728 487840 105780 487892
rect 215392 487840 215444 487892
rect 232504 487840 232556 487892
rect 299204 487840 299256 487892
rect 101128 487772 101180 487824
rect 211160 487772 211212 487824
rect 212448 487772 212500 487824
rect 232596 487772 232648 487824
rect 299296 487772 299348 487824
rect 312544 487772 312596 487824
rect 313004 487772 313056 487824
rect 408132 487772 408184 487824
rect 319628 487636 319680 487688
rect 427820 487636 427872 487688
rect 326344 487568 326396 487620
rect 434720 487568 434772 487620
rect 318064 487500 318116 487552
rect 426440 487500 426492 487552
rect 204444 487432 204496 487484
rect 222844 487432 222896 487484
rect 322940 487432 322992 487484
rect 433340 487432 433392 487484
rect 102416 487364 102468 487416
rect 211804 487364 211856 487416
rect 212448 487364 212500 487416
rect 226984 487364 227036 487416
rect 324964 487364 325016 487416
rect 434720 487364 434772 487416
rect 100024 487296 100076 487348
rect 210424 487296 210476 487348
rect 214840 487296 214892 487348
rect 229744 487296 229796 487348
rect 320916 487296 320968 487348
rect 430580 487296 430632 487348
rect 98920 487228 98972 487280
rect 209044 487228 209096 487280
rect 213736 487228 213788 487280
rect 229836 487228 229888 487280
rect 320088 487228 320140 487280
rect 429200 487228 429252 487280
rect 97816 487160 97868 487212
rect 207664 487160 207716 487212
rect 215392 487160 215444 487212
rect 244924 487160 244976 487212
rect 321560 487160 321612 487212
rect 322204 487160 322256 487212
rect 432144 487160 432196 487212
rect 457444 487160 457496 487212
rect 465080 487160 465132 487212
rect 299388 487092 299440 487144
rect 311900 487092 311952 487144
rect 312544 487092 312596 487144
rect 243544 486616 243596 486668
rect 322940 486616 322992 486668
rect 172244 486548 172296 486600
rect 254860 486548 254912 486600
rect 187700 486480 187752 486532
rect 235264 486480 235316 486532
rect 253940 486480 253992 486532
rect 409420 486480 409472 486532
rect 216772 486412 216824 486464
rect 542360 486412 542412 486464
rect 297272 486004 297324 486056
rect 297732 486004 297784 486056
rect 296812 485936 296864 485988
rect 297916 485936 297968 485988
rect 243636 485800 243688 485852
rect 244648 485800 244700 485852
rect 240784 485120 240836 485172
rect 320916 485120 320968 485172
rect 173256 485052 173308 485104
rect 247224 485052 247276 485104
rect 248420 485052 248472 485104
rect 409328 485052 409380 485104
rect 221464 484372 221516 484424
rect 580172 484372 580224 484424
rect 251640 483692 251692 483744
rect 409236 483692 409288 483744
rect 216956 483624 217008 483676
rect 580264 483624 580316 483676
rect 242164 482400 242216 482452
rect 321560 482400 321612 482452
rect 106004 482332 106056 482384
rect 234620 482332 234672 482384
rect 246396 482332 246448 482384
rect 360200 482332 360252 482384
rect 216680 482264 216732 482316
rect 501604 482264 501656 482316
rect 173164 481040 173216 481092
rect 250996 481040 251048 481092
rect 236092 480972 236144 481024
rect 434720 480972 434772 481024
rect 215300 480904 215352 480956
rect 516784 480904 516836 480956
rect 238116 479680 238168 479732
rect 319628 479680 319680 479732
rect 238852 479612 238904 479664
rect 339500 479612 339552 479664
rect 126888 479544 126940 479596
rect 240876 479544 240928 479596
rect 215484 479476 215536 479528
rect 514024 479476 514076 479528
rect 172152 478320 172204 478372
rect 248512 478320 248564 478372
rect 246488 478252 246540 478304
rect 354680 478252 354732 478304
rect 246764 478184 246816 478236
rect 406476 478184 406528 478236
rect 218244 478116 218296 478168
rect 395344 478116 395396 478168
rect 235264 477368 235316 477420
rect 293408 477436 293460 477488
rect 218152 476824 218204 476876
rect 403624 476824 403676 476876
rect 210424 476756 210476 476808
rect 239404 476756 239456 476808
rect 241612 476756 241664 476808
rect 459560 476756 459612 476808
rect 234804 476076 234856 476128
rect 235264 476076 235316 476128
rect 244372 476008 244424 476060
rect 244924 476008 244976 476060
rect 326344 476008 326396 476060
rect 236276 475396 236328 475448
rect 329840 475396 329892 475448
rect 217140 475328 217192 475380
rect 527180 475328 527232 475380
rect 3240 474716 3292 474768
rect 40684 474716 40736 474768
rect 235908 474648 235960 474700
rect 240968 474648 241020 474700
rect 241428 474648 241480 474700
rect 242256 474648 242308 474700
rect 244924 474104 244976 474156
rect 324964 474104 325016 474156
rect 77944 474036 77996 474088
rect 229928 474036 229980 474088
rect 237932 474036 237984 474088
rect 335360 474036 335412 474088
rect 215668 473968 215720 474020
rect 512644 473968 512696 474020
rect 216588 472744 216640 472796
rect 235540 472744 235592 472796
rect 236644 472744 236696 472796
rect 318064 472744 318116 472796
rect 32404 472676 32456 472728
rect 224316 472676 224368 472728
rect 238024 472676 238076 472728
rect 324320 472676 324372 472728
rect 215392 472608 215444 472660
rect 511264 472608 511316 472660
rect 211804 471928 211856 471980
rect 241704 471928 241756 471980
rect 242164 471928 242216 471980
rect 40684 471248 40736 471300
rect 224500 471248 224552 471300
rect 237472 471248 237524 471300
rect 440240 471248 440292 471300
rect 214012 470568 214064 470620
rect 579988 470568 580040 470620
rect 207664 470500 207716 470552
rect 236644 470500 236696 470552
rect 10324 469888 10376 469940
rect 224684 469888 224736 469940
rect 239036 469888 239088 469940
rect 449900 469888 449952 469940
rect 217324 469820 217376 469872
rect 509884 469820 509936 469872
rect 219624 468596 219676 468648
rect 296076 468596 296128 468648
rect 218336 468528 218388 468580
rect 399484 468528 399536 468580
rect 22744 468460 22796 468512
rect 223764 468460 223816 468512
rect 238760 468460 238812 468512
rect 444380 468460 444432 468512
rect 178684 467236 178736 467288
rect 221372 467236 221424 467288
rect 218428 467168 218480 467220
rect 409144 467168 409196 467220
rect 121368 467100 121420 467152
rect 239496 467100 239548 467152
rect 244556 467100 244608 467152
rect 470600 467100 470652 467152
rect 136548 465808 136600 465860
rect 243360 465808 243412 465860
rect 217508 465740 217560 465792
rect 406384 465740 406436 465792
rect 243084 465672 243136 465724
rect 457444 465672 457496 465724
rect 220728 464516 220780 464568
rect 237012 464516 237064 464568
rect 231492 464448 231544 464500
rect 311900 464448 311952 464500
rect 4068 464380 4120 464432
rect 224224 464380 224276 464432
rect 240324 464380 240376 464432
rect 454684 464380 454736 464432
rect 215852 464312 215904 464364
rect 504364 464312 504416 464364
rect 209044 463632 209096 463684
rect 237564 463632 237616 463684
rect 238116 463632 238168 463684
rect 219716 463156 219768 463208
rect 282920 463156 282972 463208
rect 240508 463088 240560 463140
rect 345020 463088 345072 463140
rect 230756 463020 230808 463072
rect 408224 463020 408276 463072
rect 216864 462952 216916 463004
rect 508504 462952 508556 463004
rect 2872 462340 2924 462392
rect 225604 462340 225656 462392
rect 219900 461796 219952 461848
rect 291844 461796 291896 461848
rect 131028 461728 131080 461780
rect 242072 461728 242124 461780
rect 71780 461660 71832 461712
rect 221556 461660 221608 461712
rect 241796 461660 241848 461712
rect 349160 461660 349212 461712
rect 215760 461592 215812 461644
rect 507124 461592 507176 461644
rect 239404 460776 239456 460828
rect 319444 460844 319496 460896
rect 218612 460300 218664 460352
rect 293224 460300 293276 460352
rect 14464 460232 14516 460284
rect 224040 460232 224092 460284
rect 214196 460164 214248 460216
rect 502984 460164 503036 460216
rect 203524 459484 203576 459536
rect 231584 459484 231636 459536
rect 246304 458940 246356 458992
rect 363144 458940 363196 458992
rect 171968 458872 172020 458924
rect 249800 458872 249852 458924
rect 253296 458872 253348 458924
rect 371516 458872 371568 458924
rect 40040 458804 40092 458856
rect 221004 458804 221056 458856
rect 247040 458804 247092 458856
rect 379888 458804 379940 458856
rect 299388 458736 299440 458788
rect 329656 458736 329708 458788
rect 299480 458668 299532 458720
rect 342536 458668 342588 458720
rect 296076 458600 296128 458652
rect 346400 458600 346452 458652
rect 299572 458532 299624 458584
rect 350908 458532 350960 458584
rect 298744 458464 298796 458516
rect 359280 458464 359332 458516
rect 298008 458396 298060 458448
rect 367652 458396 367704 458448
rect 355784 458328 355836 458380
rect 376024 458328 376076 458380
rect 293224 458260 293276 458312
rect 309048 458260 309100 458312
rect 299664 458192 299716 458244
rect 321284 458192 321336 458244
rect 174544 457512 174596 457564
rect 221280 457512 221332 457564
rect 6920 457444 6972 457496
rect 220820 457444 220872 457496
rect 227352 457444 227404 457496
rect 355784 457444 355836 457496
rect 222936 457240 222988 457292
rect 317420 457240 317472 457292
rect 228456 457172 228508 457224
rect 325792 457172 325844 457224
rect 236368 457104 236420 457156
rect 338028 457104 338080 457156
rect 228364 457036 228416 457088
rect 334164 457036 334216 457088
rect 247132 456968 247184 457020
rect 354772 456968 354824 457020
rect 223028 456900 223080 456952
rect 383752 456900 383804 456952
rect 223856 456764 223908 456816
rect 224316 456764 224368 456816
rect 385500 456832 385552 456884
rect 299020 456764 299072 456816
rect 580172 456764 580224 456816
rect 240508 456084 240560 456136
rect 241152 456084 241204 456136
rect 299756 456084 299808 456136
rect 300768 456084 300820 456136
rect 235080 456016 235132 456068
rect 312636 456016 312688 456068
rect 252652 455948 252704 456000
rect 385316 455948 385368 456000
rect 251732 455880 251784 455932
rect 385408 455880 385460 455932
rect 251364 455812 251416 455864
rect 385040 455812 385092 455864
rect 250168 455744 250220 455796
rect 384120 455744 384172 455796
rect 244464 455676 244516 455728
rect 384212 455676 384264 455728
rect 298928 455608 298980 455660
rect 300308 455608 300360 455660
rect 300768 455608 300820 455660
rect 385224 455608 385276 455660
rect 237748 455540 237800 455592
rect 384028 455540 384080 455592
rect 214288 455472 214340 455524
rect 384304 455472 384356 455524
rect 214472 455404 214524 455456
rect 580264 455404 580316 455456
rect 299848 455336 299900 455388
rect 304172 455336 304224 455388
rect 248696 454860 248748 454912
rect 299848 454860 299900 454912
rect 234712 454792 234764 454844
rect 299572 454792 299624 454844
rect 235264 454724 235316 454776
rect 299480 454724 299532 454776
rect 219072 454656 219124 454708
rect 295984 454656 296036 454708
rect 182824 453432 182876 453484
rect 221096 453432 221148 453484
rect 215944 453364 215996 453416
rect 284944 453364 284996 453416
rect 214656 453296 214708 453348
rect 299020 453296 299072 453348
rect 237564 453092 237616 453144
rect 237840 453092 237892 453144
rect 254124 452548 254176 452600
rect 282092 452548 282144 452600
rect 243176 452480 243228 452532
rect 247040 452480 247092 452532
rect 255872 452480 255924 452532
rect 284300 452480 284352 452532
rect 254584 452412 254636 452464
rect 284392 452412 284444 452464
rect 253204 452344 253256 452396
rect 284484 452344 284536 452396
rect 250720 452276 250772 452328
rect 283012 452276 283064 452328
rect 251548 452208 251600 452260
rect 284576 452208 284628 452260
rect 219716 452140 219768 452192
rect 219992 452140 220044 452192
rect 248144 452140 248196 452192
rect 281632 452140 281684 452192
rect 249432 452072 249484 452124
rect 283104 452072 283156 452124
rect 245844 452004 245896 452056
rect 280988 452004 281040 452056
rect 171784 451936 171836 451988
rect 220728 451936 220780 451988
rect 234620 451936 234672 451988
rect 235632 451936 235684 451988
rect 239036 451936 239088 451988
rect 240048 451936 240100 451988
rect 241612 451936 241664 451988
rect 242624 451936 242676 451988
rect 243084 451936 243136 451988
rect 243912 451936 243964 451988
rect 247408 451936 247460 451988
rect 299388 451936 299440 451988
rect 217324 451868 217376 451920
rect 286324 451868 286376 451920
rect 214840 451256 214892 451308
rect 221464 451256 221516 451308
rect 233976 451256 234028 451308
rect 297824 451256 297876 451308
rect 229836 451188 229888 451240
rect 242992 451188 243044 451240
rect 243544 451188 243596 451240
rect 189080 450916 189132 450968
rect 230848 450916 230900 450968
rect 188436 450848 188488 450900
rect 234252 450848 234304 450900
rect 187332 450780 187384 450832
rect 233792 450780 233844 450832
rect 256056 450780 256108 450832
rect 293224 450780 293276 450832
rect 187148 450712 187200 450764
rect 233424 450712 233476 450764
rect 254768 450712 254820 450764
rect 298008 450712 298060 450764
rect 187516 450644 187568 450696
rect 234068 450644 234120 450696
rect 255688 450644 255740 450696
rect 299756 450644 299808 450696
rect 187424 450576 187476 450628
rect 255320 450576 255372 450628
rect 187240 450508 187292 450560
rect 255412 450508 255464 450560
rect 3516 449828 3568 449880
rect 223028 449828 223080 449880
rect 229744 449828 229796 449880
rect 244924 449828 244976 449880
rect 204904 449760 204956 449812
rect 232596 449760 232648 449812
rect 187056 449692 187108 449744
rect 232780 449692 232832 449744
rect 238116 449692 238168 449744
rect 187608 449624 187660 449676
rect 233056 449624 233108 449676
rect 239588 449624 239640 449676
rect 190000 449556 190052 449608
rect 246120 449556 246172 449608
rect 253848 449556 253900 449608
rect 281080 449556 281132 449608
rect 189908 449488 189960 449540
rect 247316 449488 247368 449540
rect 252560 449488 252612 449540
rect 281816 449488 281868 449540
rect 171876 449420 171928 449472
rect 252376 449420 252428 449472
rect 140688 449352 140740 449404
rect 244648 449352 244700 449404
rect 251272 449352 251324 449404
rect 281908 449420 281960 449472
rect 115848 449284 115900 449336
rect 238208 449284 238260 449336
rect 249892 449284 249944 449336
rect 282000 449352 282052 449404
rect 252744 449284 252796 449336
rect 281724 449284 281776 449336
rect 111708 449216 111760 449268
rect 236920 449216 236972 449268
rect 246672 449216 246724 449268
rect 298744 449216 298796 449268
rect 3884 449148 3936 449200
rect 223120 449148 223172 449200
rect 241520 449148 241572 449200
rect 298928 449148 298980 449200
rect 248696 449080 248748 449132
rect 252744 449080 252796 449132
rect 255412 448944 255464 448996
rect 293592 448944 293644 448996
rect 252192 448876 252244 448928
rect 293684 448876 293736 448928
rect 249616 448808 249668 448860
rect 293224 448808 293276 448860
rect 244280 448740 244332 448792
rect 244924 448740 244976 448792
rect 247040 448740 247092 448792
rect 293868 448740 293920 448792
rect 244096 448672 244148 448724
rect 296536 448672 296588 448724
rect 230480 448604 230532 448656
rect 293408 448604 293460 448656
rect 230296 448536 230348 448588
rect 293776 448536 293828 448588
rect 23480 448468 23532 448520
rect 222200 448468 222252 448520
rect 222936 448468 222988 448520
rect 238116 448468 238168 448520
rect 297640 448468 297692 448520
rect 239588 448400 239640 448452
rect 297732 448400 297784 448452
rect 222844 448332 222896 448384
rect 231952 448332 232004 448384
rect 232504 448332 232556 448384
rect 233424 448264 233476 448316
rect 297916 448332 297968 448384
rect 184204 448196 184256 448248
rect 221648 448196 221700 448248
rect 226984 448196 227036 448248
rect 240416 448196 240468 448248
rect 3976 448128 4028 448180
rect 223488 448128 223540 448180
rect 233792 448128 233844 448180
rect 297456 448264 297508 448316
rect 255320 448196 255372 448248
rect 256240 448196 256292 448248
rect 297548 448196 297600 448248
rect 3700 448060 3752 448112
rect 222936 448060 222988 448112
rect 3608 447992 3660 448044
rect 222568 447992 222620 448044
rect 3792 447924 3844 447976
rect 223304 447924 223356 447976
rect 231768 447924 231820 447976
rect 239680 447924 239732 447976
rect 3424 447856 3476 447908
rect 222384 447856 222436 447908
rect 236736 447856 236788 447908
rect 253296 447856 253348 447908
rect 3240 447788 3292 447840
rect 224776 447788 224828 447840
rect 226248 447788 226300 447840
rect 238392 447788 238444 447840
rect 245752 447788 245804 447840
rect 296076 447788 296128 447840
rect 246212 447720 246264 447772
rect 246488 447720 246540 447772
rect 244740 447652 244792 447704
rect 249984 447652 250036 447704
rect 240600 447584 240652 447636
rect 230112 447516 230164 447568
rect 219440 447380 219492 447432
rect 219900 447380 219952 447432
rect 231768 447380 231820 447432
rect 214012 447312 214064 447364
rect 215024 447312 215076 447364
rect 215300 447312 215352 447364
rect 216128 447312 216180 447364
rect 217140 447312 217192 447364
rect 217600 447312 217652 447364
rect 218060 447312 218112 447364
rect 218888 447312 218940 447364
rect 221004 447312 221056 447364
rect 221832 447312 221884 447364
rect 214196 447244 214248 447296
rect 215208 447244 215260 447296
rect 215852 447244 215904 447296
rect 216312 447244 216364 447296
rect 216772 447244 216824 447296
rect 217784 447244 217836 447296
rect 218612 447244 218664 447296
rect 219256 447244 219308 447296
rect 220912 447244 220964 447296
rect 221372 447244 221424 447296
rect 224224 447244 224276 447296
rect 224684 447244 224736 447296
rect 241888 447516 241940 447568
rect 246304 447516 246356 447568
rect 244372 447448 244424 447500
rect 245568 447448 245620 447500
rect 245844 447448 245896 447500
rect 246856 447448 246908 447500
rect 251364 447516 251416 447568
rect 251824 447516 251876 447568
rect 298008 447448 298060 447500
rect 235448 447380 235500 447432
rect 293500 447380 293552 447432
rect 293132 447312 293184 447364
rect 296628 447244 296680 447296
rect 220820 447176 220872 447228
rect 222016 447176 222068 447228
rect 223304 447176 223356 447228
rect 298652 447176 298704 447228
rect 213368 447108 213420 447160
rect 296260 447108 296312 447160
rect 229928 447040 229980 447092
rect 230664 447040 230716 447092
rect 243728 447040 243780 447092
rect 246212 447040 246264 447092
rect 250352 446972 250404 447024
rect 282276 447040 282328 447092
rect 247776 446904 247828 446956
rect 258540 446904 258592 446956
rect 250168 446836 250220 446888
rect 283564 446972 283616 447024
rect 258908 446904 258960 446956
rect 282184 446904 282236 446956
rect 258816 446836 258868 446888
rect 285036 446836 285088 446888
rect 224960 446768 225012 446820
rect 225604 446768 225656 446820
rect 248972 446768 249024 446820
rect 251456 446768 251508 446820
rect 289176 446768 289228 446820
rect 4988 446700 5040 446752
rect 227720 446700 227772 446752
rect 252744 446700 252796 446752
rect 293316 446700 293368 446752
rect 4804 446632 4856 446684
rect 228824 446632 228876 446684
rect 246396 446632 246448 446684
rect 287704 446632 287756 446684
rect 3516 446564 3568 446616
rect 229376 446564 229428 446616
rect 247592 446564 247644 446616
rect 289084 446564 289136 446616
rect 188988 446496 189040 446548
rect 220544 446496 220596 446548
rect 238116 446496 238168 446548
rect 255412 446496 255464 446548
rect 256608 446496 256660 446548
rect 298100 446496 298152 446548
rect 188896 446428 188948 446480
rect 220360 446428 220412 446480
rect 233240 446428 233292 446480
rect 251732 446428 251784 446480
rect 256516 446428 256568 446480
rect 299848 446428 299900 446480
rect 172060 446360 172112 446412
rect 245936 446360 245988 446412
rect 253940 446360 253992 446412
rect 298836 446360 298888 446412
rect 3608 446292 3660 446344
rect 228640 446292 228692 446344
rect 255320 446292 255372 446344
rect 286416 446292 286468 446344
rect 209136 446224 209188 446276
rect 230388 446224 230440 446276
rect 252928 446224 252980 446276
rect 282368 446224 282420 446276
rect 221648 446156 221700 446208
rect 246948 446156 247000 446208
rect 248880 446156 248932 446208
rect 258816 446156 258868 446208
rect 5172 446088 5224 446140
rect 226064 446088 226116 446140
rect 234344 446088 234396 446140
rect 256332 446088 256384 446140
rect 5080 446020 5132 446072
rect 226616 446020 226668 446072
rect 216588 445952 216640 446004
rect 225512 445952 225564 446004
rect 213828 445884 213880 445936
rect 228088 445884 228140 445936
rect 211068 445816 211120 445868
rect 226984 445816 227036 445868
rect 232872 445816 232924 445868
rect 249892 445952 249944 446004
rect 245384 445884 245436 445936
rect 245016 445816 245068 445868
rect 246304 445816 246356 445868
rect 256516 445816 256568 445868
rect 208400 445748 208452 445800
rect 227536 445748 227588 445800
rect 236000 445748 236052 445800
rect 238024 445748 238076 445800
rect 240232 445748 240284 445800
rect 295892 445748 295944 445800
rect 227904 445680 227956 445732
rect 228456 445680 228508 445732
rect 196624 445544 196676 445596
rect 227904 445544 227956 445596
rect 225512 445476 225564 445528
rect 266176 445476 266228 445528
rect 199660 445408 199712 445460
rect 226248 445408 226300 445460
rect 196716 445340 196768 445392
rect 226800 445340 226852 445392
rect 254124 445340 254176 445392
rect 255136 445340 255188 445392
rect 210792 445272 210844 445324
rect 273904 445272 273956 445324
rect 199568 445204 199620 445256
rect 227352 445204 227404 445256
rect 236276 445204 236328 445256
rect 237288 445204 237340 445256
rect 237932 445204 237984 445256
rect 238576 445204 238628 445256
rect 238852 445204 238904 445256
rect 239864 445204 239916 445256
rect 240324 445204 240376 445256
rect 241336 445204 241388 445256
rect 241796 445204 241848 445256
rect 242440 445204 242492 445256
rect 247132 445204 247184 445256
rect 248328 445204 248380 445256
rect 248420 445204 248472 445256
rect 249064 445204 249116 445256
rect 3792 445136 3844 445188
rect 208400 445136 208452 445188
rect 213552 445136 213604 445188
rect 269856 445136 269908 445188
rect 3884 445068 3936 445120
rect 211068 445068 211120 445120
rect 215668 445068 215720 445120
rect 216496 445068 216548 445120
rect 217048 445068 217100 445120
rect 217324 445068 217376 445120
rect 218244 445068 218296 445120
rect 218704 445068 218756 445120
rect 229560 445068 229612 445120
rect 268476 445068 268528 445120
rect 3700 445000 3752 445052
rect 213828 445000 213880 445052
rect 246948 445000 247000 445052
rect 299480 445000 299532 445052
rect 226800 444932 226852 444984
rect 267096 444932 267148 444984
rect 199476 444864 199528 444916
rect 228456 444864 228508 444916
rect 212448 444796 212500 444848
rect 268384 444796 268436 444848
rect 211344 444728 211396 444780
rect 275284 444728 275336 444780
rect 210976 444660 211028 444712
rect 278044 444660 278096 444712
rect 213920 444592 213972 444644
rect 296444 444592 296496 444644
rect 213736 444524 213788 444576
rect 299296 444524 299348 444576
rect 98644 444456 98696 444508
rect 225696 444456 225748 444508
rect 253480 444456 253532 444508
rect 293316 444456 293368 444508
rect 13084 444388 13136 444440
rect 225144 444388 225196 444440
rect 254400 444388 254452 444440
rect 266084 444388 266136 444440
rect 251548 444184 251600 444236
rect 252008 444184 252060 444236
rect 213000 444048 213052 444100
rect 220268 444048 220320 444100
rect 256516 443844 256568 443896
rect 295800 443844 295852 443896
rect 214196 443776 214248 443828
rect 217508 443776 217560 443828
rect 254492 443776 254544 443828
rect 256148 443776 256200 443828
rect 256332 443776 256384 443828
rect 297364 443776 297416 443828
rect 249892 443708 249944 443760
rect 297456 443708 297508 443760
rect 3240 443640 3292 443692
rect 216588 443640 216640 443692
rect 212540 443572 212592 443624
rect 229836 443640 229888 443692
rect 234436 443640 234488 443692
rect 239956 443640 240008 443692
rect 199384 443436 199436 443488
rect 212540 443436 212592 443488
rect 4068 443232 4120 443284
rect 3332 443164 3384 443216
rect 215852 443368 215904 443420
rect 220268 443504 220320 443556
rect 216588 443368 216640 443420
rect 217508 443368 217560 443420
rect 234436 443436 234488 443488
rect 239036 443504 239088 443556
rect 242716 443640 242768 443692
rect 248972 443640 249024 443692
rect 297548 443640 297600 443692
rect 242900 443504 242952 443556
rect 225236 443368 225288 443420
rect 225788 443368 225840 443420
rect 226340 443368 226392 443420
rect 228180 443368 228232 443420
rect 3976 443096 4028 443148
rect 4896 443028 4948 443080
rect 3424 442960 3476 443012
rect 229468 443368 229520 443420
rect 233700 443368 233752 443420
rect 239220 443368 239272 443420
rect 239956 443368 240008 443420
rect 242716 443368 242768 443420
rect 254492 443368 254544 443420
rect 256148 443368 256200 443420
rect 265992 443368 266044 443420
rect 298560 443300 298612 443352
rect 266360 443232 266412 443284
rect 265532 443096 265584 443148
rect 267004 443028 267056 443080
rect 298008 442960 298060 443012
rect 266360 440172 266412 440224
rect 298008 440172 298060 440224
rect 265532 436024 265584 436076
rect 297180 436024 297232 436076
rect 267096 431876 267148 431928
rect 298008 431876 298060 431928
rect 384304 431876 384356 431928
rect 580172 431876 580224 431928
rect 268476 426368 268528 426420
rect 298008 426368 298060 426420
rect 3148 423580 3200 423632
rect 13084 423580 13136 423632
rect 267004 408416 267056 408468
rect 298008 408416 298060 408468
rect 266176 404268 266228 404320
rect 298008 404268 298060 404320
rect 299572 401208 299624 401260
rect 293868 401072 293920 401124
rect 299664 401072 299716 401124
rect 293776 401004 293828 401056
rect 299480 401004 299532 401056
rect 293592 400936 293644 400988
rect 299572 400936 299624 400988
rect 293684 400868 293736 400920
rect 299572 400732 299624 400784
rect 299848 400732 299900 400784
rect 299480 400664 299532 400716
rect 299664 400596 299716 400648
rect 307576 400596 307628 400648
rect 311900 400596 311952 400648
rect 324228 400596 324280 400648
rect 340972 400596 341024 400648
rect 298560 400120 298612 400172
rect 579988 400120 580040 400172
rect 293316 400052 293368 400104
rect 385040 400052 385092 400104
rect 217232 399168 217284 399220
rect 216956 399032 217008 399084
rect 217232 399032 217284 399084
rect 244372 399100 244424 399152
rect 437480 399100 437532 399152
rect 217600 398964 217652 399016
rect 208032 398760 208084 398812
rect 210056 398760 210108 398812
rect 210240 398760 210292 398812
rect 207664 398692 207716 398744
rect 207940 398624 207992 398676
rect 210148 398624 210200 398676
rect 214012 398624 214064 398676
rect 214472 398624 214524 398676
rect 207020 398556 207072 398608
rect 207848 398488 207900 398540
rect 210240 398488 210292 398540
rect 203524 398420 203576 398472
rect 211804 398420 211856 398472
rect 209228 398352 209280 398404
rect 212172 398352 212224 398404
rect 217692 398896 217744 398948
rect 217508 398692 217560 398744
rect 217600 398692 217652 398744
rect 219348 398964 219400 399016
rect 219440 398964 219492 399016
rect 236092 398896 236144 398948
rect 253664 399032 253716 399084
rect 277400 399032 277452 399084
rect 256056 398964 256108 399016
rect 299480 398964 299532 399016
rect 230848 398760 230900 398812
rect 331220 398896 331272 398948
rect 217232 398624 217284 398676
rect 217784 398624 217836 398676
rect 229284 398624 229336 398676
rect 230020 398624 230072 398676
rect 244832 398692 244884 398744
rect 263600 398828 263652 398880
rect 296628 398760 296680 398812
rect 379244 398760 379296 398812
rect 217784 398488 217836 398540
rect 222844 398488 222896 398540
rect 228456 398488 228508 398540
rect 230020 398488 230072 398540
rect 233608 398488 233660 398540
rect 239864 398556 239916 398608
rect 245660 398556 245712 398608
rect 256056 398692 256108 398744
rect 295892 398692 295944 398744
rect 303896 398692 303948 398744
rect 255504 398624 255556 398676
rect 269764 398624 269816 398676
rect 299572 398624 299624 398676
rect 374736 398624 374788 398676
rect 261484 398556 261536 398608
rect 293224 398556 293276 398608
rect 366364 398556 366416 398608
rect 245936 398488 245988 398540
rect 264244 398488 264296 398540
rect 299388 398488 299440 398540
rect 370872 398488 370924 398540
rect 223396 398420 223448 398472
rect 233332 398420 233384 398472
rect 239864 398420 239916 398472
rect 240416 398420 240468 398472
rect 245384 398420 245436 398472
rect 246212 398420 246264 398472
rect 264336 398420 264388 398472
rect 296536 398420 296588 398472
rect 362500 398420 362552 398472
rect 226432 398352 226484 398404
rect 204904 398284 204956 398336
rect 212264 398284 212316 398336
rect 213368 398284 213420 398336
rect 223120 398284 223172 398336
rect 229744 398284 229796 398336
rect 241520 398284 241572 398336
rect 249064 398284 249116 398336
rect 252652 398284 252704 398336
rect 171140 398216 171192 398268
rect 223672 398216 223724 398268
rect 230572 398216 230624 398268
rect 125600 398148 125652 398200
rect 220084 398148 220136 398200
rect 242072 398148 242124 398200
rect 24860 398080 24912 398132
rect 204904 398080 204956 398132
rect 209780 398080 209832 398132
rect 210700 398080 210752 398132
rect 212448 398080 212500 398132
rect 225052 398080 225104 398132
rect 210148 398012 210200 398064
rect 218336 398012 218388 398064
rect 210056 397944 210108 397996
rect 218888 397944 218940 397996
rect 238208 397944 238260 397996
rect 211528 397876 211580 397928
rect 217232 397876 217284 397928
rect 219440 397876 219492 397928
rect 239312 397944 239364 397996
rect 242624 397944 242676 397996
rect 245660 398080 245712 398132
rect 246488 398080 246540 398132
rect 247684 398080 247736 398132
rect 247960 398080 248012 398132
rect 244280 398012 244332 398064
rect 255596 398352 255648 398404
rect 275376 398352 275428 398404
rect 295800 398352 295852 398404
rect 357992 398352 358044 398404
rect 257528 398284 257580 398336
rect 264980 398284 265032 398336
rect 293500 398284 293552 398336
rect 349620 398284 349672 398336
rect 256700 398216 256752 398268
rect 298652 398216 298704 398268
rect 329012 398216 329064 398268
rect 543740 398148 543792 398200
rect 254308 398080 254360 398132
rect 564440 398080 564492 398132
rect 259552 398012 259604 398064
rect 293408 398012 293460 398064
rect 320640 398012 320692 398064
rect 206284 397808 206336 397860
rect 236368 397808 236420 397860
rect 239312 397808 239364 397860
rect 210240 397740 210292 397792
rect 216956 397740 217008 397792
rect 217048 397740 217100 397792
rect 217784 397740 217836 397792
rect 219440 397740 219492 397792
rect 227444 397740 227496 397792
rect 193220 397672 193272 397724
rect 225328 397672 225380 397724
rect 228272 397672 228324 397724
rect 230480 397672 230532 397724
rect 231952 397672 232004 397724
rect 244832 397876 244884 397928
rect 245936 397876 245988 397928
rect 243176 397808 243228 397860
rect 258816 397944 258868 397996
rect 266084 397944 266136 397996
rect 316132 397944 316184 397996
rect 264980 397876 265032 397928
rect 345756 397876 345808 397928
rect 243728 397740 243780 397792
rect 256424 397808 256476 397860
rect 217784 397604 217836 397656
rect 220820 397604 220872 397656
rect 222200 397604 222252 397656
rect 227628 397604 227680 397656
rect 234068 397604 234120 397656
rect 244832 397672 244884 397724
rect 244464 397604 244516 397656
rect 256608 397740 256660 397792
rect 245936 397672 245988 397724
rect 246764 397672 246816 397724
rect 249064 397672 249116 397724
rect 256516 397672 256568 397724
rect 257620 397604 257672 397656
rect 209044 397536 209096 397588
rect 210792 397536 210844 397588
rect 210240 397468 210292 397520
rect 210700 397468 210752 397520
rect 211528 397536 211580 397588
rect 211896 397536 211948 397588
rect 215024 397536 215076 397588
rect 211160 397468 211212 397520
rect 213552 397468 213604 397520
rect 210792 397400 210844 397452
rect 215024 397400 215076 397452
rect 218796 397536 218848 397588
rect 218888 397536 218940 397588
rect 220728 397536 220780 397588
rect 224960 397536 225012 397588
rect 227168 397536 227220 397588
rect 239312 397536 239364 397588
rect 240048 397536 240100 397588
rect 220084 397468 220136 397520
rect 222384 397468 222436 397520
rect 225052 397468 225104 397520
rect 225604 397468 225656 397520
rect 226432 397468 226484 397520
rect 227720 397468 227772 397520
rect 231492 397468 231544 397520
rect 234068 397468 234120 397520
rect 234344 397468 234396 397520
rect 238760 397468 238812 397520
rect 240968 397468 241020 397520
rect 242624 397468 242676 397520
rect 248788 397536 248840 397588
rect 244004 397468 244056 397520
rect 244464 397468 244516 397520
rect 253664 397468 253716 397520
rect 217232 397400 217284 397452
rect 226616 397400 226668 397452
rect 257436 397536 257488 397588
rect 254032 397468 254084 397520
rect 256332 397468 256384 397520
rect 211620 397332 211672 397384
rect 218612 397332 218664 397384
rect 201500 397264 201552 397316
rect 226064 397332 226116 397384
rect 212540 397196 212592 397248
rect 213460 397196 213512 397248
rect 194600 397128 194652 397180
rect 225512 397264 225564 397316
rect 247040 397196 247092 397248
rect 247592 397196 247644 397248
rect 247684 397196 247736 397248
rect 256148 397196 256200 397248
rect 227812 397128 227864 397180
rect 229008 397128 229060 397180
rect 235448 397128 235500 397180
rect 235632 397128 235684 397180
rect 238760 397128 238812 397180
rect 239404 397128 239456 397180
rect 241704 397128 241756 397180
rect 249064 397128 249116 397180
rect 160100 397060 160152 397112
rect 222752 397060 222804 397112
rect 246212 397060 246264 397112
rect 256056 397128 256108 397180
rect 144920 396992 144972 397044
rect 221648 396992 221700 397044
rect 227812 396992 227864 397044
rect 228732 396992 228784 397044
rect 231860 396992 231912 397044
rect 232872 396992 232924 397044
rect 234896 396992 234948 397044
rect 235448 396992 235500 397044
rect 238852 396992 238904 397044
rect 239404 396992 239456 397044
rect 135260 396924 135312 396976
rect 217784 396924 217836 396976
rect 229744 396924 229796 396976
rect 131120 396856 131172 396908
rect 220544 396856 220596 396908
rect 228088 396856 228140 396908
rect 228732 396856 228784 396908
rect 230572 396856 230624 396908
rect 231584 396856 231636 396908
rect 231860 396856 231912 396908
rect 232504 396856 232556 396908
rect 233332 396856 233384 396908
rect 233700 396856 233752 396908
rect 106280 396788 106332 396840
rect 211620 396788 211672 396840
rect 212724 396788 212776 396840
rect 213184 396788 213236 396840
rect 229376 396788 229428 396840
rect 230112 396788 230164 396840
rect 231952 396788 232004 396840
rect 232320 396788 232372 396840
rect 237380 396924 237432 396976
rect 238392 396924 238444 396976
rect 238944 396924 238996 396976
rect 239312 396924 239364 396976
rect 240784 396924 240836 396976
rect 241428 396924 241480 396976
rect 234620 396856 234672 396908
rect 234988 396856 235040 396908
rect 237012 396856 237064 396908
rect 242256 396856 242308 396908
rect 242440 396788 242492 396840
rect 242808 396788 242860 396840
rect 243544 396788 243596 396840
rect 342260 396856 342312 396908
rect 40040 396720 40092 396772
rect 212540 396720 212592 396772
rect 212908 396720 212960 396772
rect 213368 396720 213420 396772
rect 214104 396720 214156 396772
rect 214564 396720 214616 396772
rect 226708 396720 226760 396772
rect 227168 396720 227220 396772
rect 229560 396720 229612 396772
rect 231032 396720 231084 396772
rect 231492 396720 231544 396772
rect 232228 396720 232280 396772
rect 209872 396652 209924 396704
rect 210516 396652 210568 396704
rect 211344 396652 211396 396704
rect 212080 396652 212132 396704
rect 212816 396652 212868 396704
rect 213828 396652 213880 396704
rect 214196 396652 214248 396704
rect 214932 396652 214984 396704
rect 225788 396652 225840 396704
rect 226248 396652 226300 396704
rect 227904 396652 227956 396704
rect 228180 396652 228232 396704
rect 228272 396652 228324 396704
rect 228824 396652 228876 396704
rect 209964 396584 210016 396636
rect 210884 396584 210936 396636
rect 211252 396584 211304 396636
rect 211988 396584 212040 396636
rect 212908 396584 212960 396636
rect 213276 396584 213328 396636
rect 214472 396584 214524 396636
rect 214748 396584 214800 396636
rect 211528 396516 211580 396568
rect 212356 396516 212408 396568
rect 213000 396516 213052 396568
rect 213644 396516 213696 396568
rect 214564 396516 214616 396568
rect 215208 396516 215260 396568
rect 226708 396516 226760 396568
rect 227260 396516 227312 396568
rect 227904 396516 227956 396568
rect 228088 396516 228140 396568
rect 229376 396516 229428 396568
rect 232688 396720 232740 396772
rect 234988 396720 235040 396772
rect 235172 396720 235224 396772
rect 235264 396720 235316 396772
rect 235908 396720 235960 396772
rect 236276 396720 236328 396772
rect 237012 396720 237064 396772
rect 237380 396720 237432 396772
rect 237748 396720 237800 396772
rect 238024 396720 238076 396772
rect 240324 396720 240376 396772
rect 240600 396720 240652 396772
rect 240784 396720 240836 396772
rect 241520 396720 241572 396772
rect 241888 396720 241940 396772
rect 243084 396720 243136 396772
rect 243360 396720 243412 396772
rect 243728 396720 243780 396772
rect 249064 396788 249116 396840
rect 402980 396788 403032 396840
rect 409880 396720 409932 396772
rect 232228 396516 232280 396568
rect 232412 396516 232464 396568
rect 232596 396516 232648 396568
rect 212632 396448 212684 396500
rect 213736 396448 213788 396500
rect 226800 396448 226852 396500
rect 227536 396448 227588 396500
rect 229468 396448 229520 396500
rect 229928 396448 229980 396500
rect 210240 396380 210292 396432
rect 210976 396380 211028 396432
rect 228088 396380 228140 396432
rect 228640 396380 228692 396432
rect 229100 396380 229152 396432
rect 229652 396380 229704 396432
rect 230848 396380 230900 396432
rect 231216 396380 231268 396432
rect 232412 396380 232464 396432
rect 236368 396652 236420 396704
rect 236736 396652 236788 396704
rect 233516 396516 233568 396568
rect 233976 396516 234028 396568
rect 234528 396516 234580 396568
rect 235080 396516 235132 396568
rect 237656 396516 237708 396568
rect 239128 396652 239180 396704
rect 239496 396652 239548 396704
rect 239036 396516 239088 396568
rect 239588 396516 239640 396568
rect 240692 396516 240744 396568
rect 243452 396516 243504 396568
rect 234804 396448 234856 396500
rect 235540 396448 235592 396500
rect 237932 396448 237984 396500
rect 238116 396448 238168 396500
rect 240140 396448 240192 396500
rect 240416 396448 240468 396500
rect 240508 396448 240560 396500
rect 241152 396448 241204 396500
rect 242900 396448 242952 396500
rect 243268 396448 243320 396500
rect 233332 396380 233384 396432
rect 233884 396380 233936 396432
rect 236092 396380 236144 396432
rect 236644 396380 236696 396432
rect 237840 396380 237892 396432
rect 238208 396380 238260 396432
rect 240324 396380 240376 396432
rect 241060 396380 241112 396432
rect 241704 396380 241756 396432
rect 241980 396380 242032 396432
rect 243176 396380 243228 396432
rect 243820 396380 243872 396432
rect 210332 396312 210384 396364
rect 211068 396312 211120 396364
rect 222752 396312 222804 396364
rect 227352 396312 227404 396364
rect 230940 396312 230992 396364
rect 231400 396312 231452 396364
rect 233240 396312 233292 396364
rect 233976 396312 234028 396364
rect 236000 396312 236052 396364
rect 236920 396312 236972 396364
rect 237564 396312 237616 396364
rect 237932 396312 237984 396364
rect 240416 396312 240468 396364
rect 241244 396312 241296 396364
rect 241612 396312 241664 396364
rect 242164 396312 242216 396364
rect 233884 396244 233936 396296
rect 234068 396244 234120 396296
rect 233240 396176 233292 396228
rect 234160 396176 234212 396228
rect 210516 396108 210568 396160
rect 217232 396108 217284 396160
rect 237656 396108 237708 396160
rect 238300 396108 238352 396160
rect 244188 396108 244240 396160
rect 245476 396108 245528 396160
rect 250444 395972 250496 396024
rect 250812 395972 250864 396024
rect 213184 395904 213236 395956
rect 213460 395904 213512 395956
rect 214012 395904 214064 395956
rect 214380 395904 214432 395956
rect 231584 395904 231636 395956
rect 256240 395904 256292 395956
rect 231492 395836 231544 395888
rect 266360 395836 266412 395888
rect 214012 395768 214064 395820
rect 214840 395768 214892 395820
rect 231308 395768 231360 395820
rect 269120 395768 269172 395820
rect 232872 395700 232924 395752
rect 276020 395700 276072 395752
rect 141424 395632 141476 395684
rect 217508 395632 217560 395684
rect 240048 395632 240100 395684
rect 333980 395632 334032 395684
rect 115940 395564 115992 395616
rect 219348 395564 219400 395616
rect 247316 395564 247368 395616
rect 247684 395564 247736 395616
rect 250168 395564 250220 395616
rect 250444 395564 250496 395616
rect 252008 395564 252060 395616
rect 535460 395564 535512 395616
rect 77300 395496 77352 395548
rect 216404 395496 216456 395548
rect 253112 395496 253164 395548
rect 549260 395496 549312 395548
rect 52460 395428 52512 395480
rect 214380 395428 214432 395480
rect 253940 395428 253992 395480
rect 560300 395428 560352 395480
rect 30380 395360 30432 395412
rect 212540 395360 212592 395412
rect 254216 395360 254268 395412
rect 564532 395360 564584 395412
rect 27620 395292 27672 395344
rect 212172 395292 212224 395344
rect 226524 395292 226576 395344
rect 226892 395292 226944 395344
rect 254768 395292 254820 395344
rect 571340 395292 571392 395344
rect 214380 395156 214432 395208
rect 214656 395156 214708 395208
rect 251548 395020 251600 395072
rect 252008 395020 252060 395072
rect 216404 394680 216456 394732
rect 223304 394680 223356 394732
rect 228364 394680 228416 394732
rect 231124 394680 231176 394732
rect 254032 394680 254084 394732
rect 254400 394680 254452 394732
rect 215300 394612 215352 394664
rect 218888 394612 218940 394664
rect 225604 394612 225656 394664
rect 227076 394612 227128 394664
rect 244556 394612 244608 394664
rect 245568 394612 245620 394664
rect 247960 394612 248012 394664
rect 258724 394612 258776 394664
rect 215392 394544 215444 394596
rect 215944 394544 215996 394596
rect 251272 394544 251324 394596
rect 251824 394544 251876 394596
rect 253940 394544 253992 394596
rect 254584 394544 254636 394596
rect 4160 394408 4212 394460
rect 209780 394408 209832 394460
rect 209136 394340 209188 394392
rect 224500 394476 224552 394528
rect 234344 394476 234396 394528
rect 305000 394476 305052 394528
rect 235632 394408 235684 394460
rect 322940 394408 322992 394460
rect 189080 394272 189132 394324
rect 212448 394272 212500 394324
rect 178040 394204 178092 394256
rect 224224 394340 224276 394392
rect 237012 394340 237064 394392
rect 332600 394340 332652 394392
rect 221096 394272 221148 394324
rect 221556 394272 221608 394324
rect 223764 394272 223816 394324
rect 224316 394272 224368 394324
rect 236828 394272 236880 394324
rect 340880 394272 340932 394324
rect 133880 394136 133932 394188
rect 215300 394136 215352 394188
rect 129740 394068 129792 394120
rect 220452 394204 220504 394256
rect 238392 394204 238444 394256
rect 347780 394204 347832 394256
rect 215576 394136 215628 394188
rect 216220 394136 216272 394188
rect 216956 394136 217008 394188
rect 217416 394136 217468 394188
rect 220912 394136 220964 394188
rect 222016 394136 222068 394188
rect 222384 394136 222436 394188
rect 222936 394136 222988 394188
rect 223856 394136 223908 394188
rect 224592 394136 224644 394188
rect 244004 394136 244056 394188
rect 365720 394136 365772 394188
rect 92480 394000 92532 394052
rect 217692 394068 217744 394120
rect 218244 394068 218296 394120
rect 218980 394068 219032 394120
rect 219532 394068 219584 394120
rect 220360 394068 220412 394120
rect 221188 394068 221240 394120
rect 221832 394068 221884 394120
rect 223948 394068 224000 394120
rect 224868 394068 224920 394120
rect 240232 394068 240284 394120
rect 382280 394068 382332 394120
rect 215668 394000 215720 394052
rect 216220 394000 216272 394052
rect 216864 394000 216916 394052
rect 217876 394000 217928 394052
rect 218612 394000 218664 394052
rect 219072 394000 219124 394052
rect 219808 394000 219860 394052
rect 220268 394000 220320 394052
rect 221556 394000 221608 394052
rect 221924 394000 221976 394052
rect 224316 394000 224368 394052
rect 224776 394000 224828 394052
rect 210424 393932 210476 393984
rect 225052 394000 225104 394052
rect 244924 394000 244976 394052
rect 252744 394000 252796 394052
rect 253112 394000 253164 394052
rect 209780 393864 209832 393916
rect 210516 393864 210568 393916
rect 215668 393864 215720 393916
rect 216312 393864 216364 393916
rect 218428 393864 218480 393916
rect 218796 393864 218848 393916
rect 219716 393864 219768 393916
rect 220176 393864 220228 393916
rect 221372 393864 221424 393916
rect 221740 393864 221792 393916
rect 222476 393864 222528 393916
rect 222936 393864 222988 393916
rect 224040 393864 224092 393916
rect 224408 393864 224460 393916
rect 216036 393796 216088 393848
rect 216588 393796 216640 393848
rect 218336 393796 218388 393848
rect 219256 393796 219308 393848
rect 219624 393796 219676 393848
rect 220636 393796 220688 393848
rect 221004 393796 221056 393848
rect 222108 393796 222160 393848
rect 244464 393796 244516 393848
rect 246304 393932 246356 393984
rect 246948 393932 247000 393984
rect 251364 393932 251416 393984
rect 251548 393932 251600 393984
rect 245568 393864 245620 393916
rect 440240 394000 440292 394052
rect 245844 393796 245896 393848
rect 246580 393796 246632 393848
rect 250076 393796 250128 393848
rect 250260 393796 250312 393848
rect 251180 393796 251232 393848
rect 251364 393796 251416 393848
rect 251640 393796 251692 393848
rect 251916 393796 251968 393848
rect 252836 393796 252888 393848
rect 253204 393796 253256 393848
rect 215484 393728 215536 393780
rect 216496 393728 216548 393780
rect 218428 393728 218480 393780
rect 219164 393728 219216 393780
rect 244372 393728 244424 393780
rect 245200 393728 245252 393780
rect 247224 393728 247276 393780
rect 215944 393660 215996 393712
rect 216404 393660 216456 393712
rect 252744 393728 252796 393780
rect 253480 393728 253532 393780
rect 251180 393660 251232 393712
rect 252100 393660 252152 393712
rect 252652 393660 252704 393712
rect 252928 393660 252980 393712
rect 248696 393592 248748 393644
rect 492680 393932 492732 393984
rect 254124 393864 254176 393916
rect 254860 393864 254912 393916
rect 247316 393524 247368 393576
rect 252928 393252 252980 393304
rect 253388 393252 253440 393304
rect 244740 393116 244792 393168
rect 245108 393116 245160 393168
rect 244648 393048 244700 393100
rect 245292 393048 245344 393100
rect 247684 393048 247736 393100
rect 253664 393048 253716 393100
rect 252560 392980 252612 393032
rect 253204 392980 253256 393032
rect 231032 392912 231084 392964
rect 267740 392912 267792 392964
rect 239588 392844 239640 392896
rect 295340 392844 295392 392896
rect 241796 392776 241848 392828
rect 401600 392776 401652 392828
rect 202880 392708 202932 392760
rect 225880 392708 225932 392760
rect 252560 392708 252612 392760
rect 253572 392708 253624 392760
rect 253664 392708 253716 392760
rect 483020 392708 483072 392760
rect 160192 392640 160244 392692
rect 217048 392640 217100 392692
rect 248512 392640 248564 392692
rect 498200 392640 498252 392692
rect 109040 392572 109092 392624
rect 214656 392572 214708 392624
rect 250444 392572 250496 392624
rect 512000 392572 512052 392624
rect 245660 392368 245712 392420
rect 246028 392368 246080 392420
rect 217140 392164 217192 392216
rect 217968 392164 218020 392216
rect 248788 392164 248840 392216
rect 249432 392164 249484 392216
rect 249984 392164 250036 392216
rect 250536 392164 250588 392216
rect 247776 392096 247828 392148
rect 224224 392028 224276 392080
rect 224684 392028 224736 392080
rect 247132 392028 247184 392080
rect 247500 392028 247552 392080
rect 247868 392028 247920 392080
rect 248420 392028 248472 392080
rect 248972 392028 249024 392080
rect 225236 391960 225288 392012
rect 229008 391960 229060 392012
rect 248420 391892 248472 391944
rect 249340 391892 249392 391944
rect 248696 391688 248748 391740
rect 249156 391688 249208 391740
rect 233424 391416 233476 391468
rect 299572 391416 299624 391468
rect 239404 391348 239456 391400
rect 365812 391348 365864 391400
rect 250812 391280 250864 391332
rect 514760 391280 514812 391332
rect 229744 391212 229796 391264
rect 250444 391212 250496 391264
rect 252008 391212 252060 391264
rect 529940 391212 529992 391264
rect 245752 391144 245804 391196
rect 246212 391144 246264 391196
rect 222752 391008 222804 391060
rect 223028 391008 223080 391060
rect 233976 389988 234028 390040
rect 293960 389988 294012 390040
rect 230020 389920 230072 389972
rect 233424 389920 233476 389972
rect 235356 389920 235408 389972
rect 316040 389920 316092 389972
rect 246764 389852 246816 389904
rect 357440 389852 357492 389904
rect 245476 389784 245528 389836
rect 438860 389784 438912 389836
rect 249800 389716 249852 389768
rect 250168 389716 250220 389768
rect 249800 389580 249852 389632
rect 250720 389580 250772 389632
rect 254308 389376 254360 389428
rect 254676 389376 254728 389428
rect 222568 389308 222620 389360
rect 223488 389308 223540 389360
rect 217324 389240 217376 389292
rect 217508 389036 217560 389088
rect 299296 379448 299348 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 98644 372512 98696 372564
rect 296444 365644 296496 365696
rect 580172 365644 580224 365696
rect 2780 358436 2832 358488
rect 5172 358436 5224 358488
rect 250352 356804 250404 356856
rect 514852 356804 514904 356856
rect 250536 356736 250588 356788
rect 517520 356736 517572 356788
rect 251824 356668 251876 356720
rect 531320 356668 531372 356720
rect 232596 355580 232648 355632
rect 281540 355580 281592 355632
rect 232504 355512 232556 355564
rect 288440 355512 288492 355564
rect 184940 355444 184992 355496
rect 224224 355444 224276 355496
rect 250168 355444 250220 355496
rect 506480 355444 506532 355496
rect 110420 355376 110472 355428
rect 208032 355376 208084 355428
rect 250260 355376 250312 355428
rect 510620 355376 510672 355428
rect 104900 355308 104952 355360
rect 218520 355308 218572 355360
rect 253296 355308 253348 355360
rect 550640 355308 550692 355360
rect 200120 354560 200172 354612
rect 225420 354560 225472 354612
rect 180800 354492 180852 354544
rect 224132 354492 224184 354544
rect 176660 354424 176712 354476
rect 224040 354424 224092 354476
rect 98000 354356 98052 354408
rect 217140 354356 217192 354408
rect 91100 354288 91152 354340
rect 216956 354288 217008 354340
rect 238116 354288 238168 354340
rect 353300 354288 353352 354340
rect 86960 354220 87012 354272
rect 217048 354220 217100 354272
rect 240876 354220 240928 354272
rect 391940 354220 391992 354272
rect 70400 354152 70452 354204
rect 212080 354152 212132 354204
rect 241980 354152 242032 354204
rect 411260 354152 411312 354204
rect 62120 354084 62172 354136
rect 214564 354084 214616 354136
rect 244832 354084 244884 354136
rect 445760 354084 445812 354136
rect 42800 354016 42852 354068
rect 213000 354016 213052 354068
rect 253204 354016 253256 354068
rect 542360 354016 542412 354068
rect 35900 353948 35952 354000
rect 213092 353948 213144 354000
rect 229652 353948 229704 354000
rect 241796 353948 241848 354000
rect 253112 353948 253164 354000
rect 546500 353948 546552 354000
rect 269856 353200 269908 353252
rect 580172 353200 580224 353252
rect 230940 352860 230992 352912
rect 270500 352860 270552 352912
rect 235172 352792 235224 352844
rect 317420 352792 317472 352844
rect 235264 352724 235316 352776
rect 321560 352724 321612 352776
rect 239312 352656 239364 352708
rect 367100 352656 367152 352708
rect 149060 352588 149112 352640
rect 221556 352588 221608 352640
rect 246580 352588 246632 352640
rect 379520 352588 379572 352640
rect 88340 352520 88392 352572
rect 210608 352520 210660 352572
rect 241888 352520 241940 352572
rect 404360 352520 404412 352572
rect 220820 351908 220872 351960
rect 226800 351908 226852 351960
rect 233792 351296 233844 351348
rect 300860 351296 300912 351348
rect 142160 351228 142212 351280
rect 221464 351228 221516 351280
rect 242624 351228 242676 351280
rect 393320 351228 393372 351280
rect 74540 351160 74592 351212
rect 216128 351160 216180 351212
rect 218520 351160 218572 351212
rect 226708 351160 226760 351212
rect 243636 351160 243688 351212
rect 423680 351160 423732 351212
rect 254492 348372 254544 348424
rect 572720 348372 572772 348424
rect 23480 338716 23532 338768
rect 209228 338716 209280 338768
rect 260104 335996 260156 336048
rect 449900 335996 449952 336048
rect 257620 334568 257672 334620
rect 429200 334568 429252 334620
rect 299112 325592 299164 325644
rect 580172 325592 580224 325644
rect 3332 320084 3384 320136
rect 199660 320084 199712 320136
rect 296260 313216 296312 313268
rect 580172 313216 580224 313268
rect 2780 306212 2832 306264
rect 5080 306212 5132 306264
rect 258816 305600 258868 305652
rect 436100 305600 436152 305652
rect 265992 299412 266044 299464
rect 580172 299412 580224 299464
rect 299204 273164 299256 273216
rect 580172 273164 580224 273216
rect 3148 267656 3200 267708
rect 196716 267656 196768 267708
rect 296352 259360 296404 259412
rect 580172 259360 580224 259412
rect 268384 245556 268436 245608
rect 580172 245556 580224 245608
rect 298928 233180 298980 233232
rect 579988 233180 580040 233232
rect 296168 219376 296220 219428
rect 580172 219376 580224 219428
rect 3056 215228 3108 215280
rect 199568 215228 199620 215280
rect 299020 206932 299072 206984
rect 579804 206932 579856 206984
rect 2780 202648 2832 202700
rect 4988 202648 5040 202700
rect 298836 193128 298888 193180
rect 580172 193128 580224 193180
rect 275376 191088 275428 191140
rect 582380 191088 582432 191140
rect 264336 188300 264388 188352
rect 460940 188300 460992 188352
rect 261484 186940 261536 186992
rect 443000 186940 443052 186992
rect 38660 180072 38712 180124
rect 202144 180072 202196 180124
rect 295984 179324 296036 179376
rect 580172 179324 580224 179376
rect 102232 178644 102284 178696
rect 207940 178644 207992 178696
rect 240784 178644 240836 178696
rect 389180 178644 389232 178696
rect 155960 177556 156012 177608
rect 222936 177556 222988 177608
rect 124220 177488 124272 177540
rect 219992 177488 220044 177540
rect 111800 177420 111852 177472
rect 218612 177420 218664 177472
rect 80060 177352 80112 177404
rect 216036 177352 216088 177404
rect 228272 177352 228324 177404
rect 232504 177352 232556 177404
rect 9680 177284 9732 177336
rect 210332 177284 210384 177336
rect 228364 177284 228416 177336
rect 235172 177284 235224 177336
rect 242256 177284 242308 177336
rect 372620 177284 372672 177336
rect 31760 168988 31812 169040
rect 203616 168988 203668 169040
rect 269764 167628 269816 167680
rect 581092 167628 581144 167680
rect 275284 166948 275336 167000
rect 580172 166948 580224 167000
rect 3056 164160 3108 164212
rect 196624 164160 196676 164212
rect 278044 153144 278096 153196
rect 580172 153144 580224 153196
rect 2780 149880 2832 149932
rect 4896 149880 4948 149932
rect 265900 139340 265952 139392
rect 580172 139340 580224 139392
rect 273904 126896 273956 126948
rect 580172 126896 580224 126948
rect 298744 113092 298796 113144
rect 579804 113092 579856 113144
rect 3332 111732 3384 111784
rect 199476 111732 199528 111784
rect 296076 100648 296128 100700
rect 580172 100648 580224 100700
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 216956 88952 217008 89004
rect 224960 88952 225012 89004
rect 232412 87728 232464 87780
rect 287060 87728 287112 87780
rect 243544 87660 243596 87712
rect 427820 87660 427872 87712
rect 251732 87592 251784 87644
rect 531412 87592 531464 87644
rect 265808 86912 265860 86964
rect 580172 86912 580224 86964
rect 240692 86300 240744 86352
rect 385040 86300 385092 86352
rect 117320 86232 117372 86284
rect 206284 86232 206336 86284
rect 246212 86232 246264 86284
rect 454040 86232 454092 86284
rect 238024 84804 238076 84856
rect 354680 84804 354732 84856
rect 233700 83580 233752 83632
rect 298100 83580 298152 83632
rect 256608 83512 256660 83564
rect 422300 83512 422352 83564
rect 243452 83444 243504 83496
rect 420920 83444 420972 83496
rect 95240 82084 95292 82136
rect 207848 82084 207900 82136
rect 249064 82084 249116 82136
rect 499580 82084 499632 82136
rect 236552 80656 236604 80708
rect 336740 80656 336792 80708
rect 265716 73108 265768 73160
rect 580172 73108 580224 73160
rect 3332 71680 3384 71732
rect 257528 71680 257580 71732
rect 283564 60664 283616 60716
rect 580172 60664 580224 60716
rect 265624 46860 265676 46912
rect 580172 46860 580224 46912
rect 162860 46248 162912 46300
rect 222752 46248 222804 46300
rect 146300 46180 146352 46232
rect 221372 46180 221424 46232
rect 229560 46180 229612 46232
rect 249064 46180 249116 46232
rect 271144 31016 271196 31068
rect 474740 31016 474792 31068
rect 264244 29588 264296 29640
rect 456800 29588 456852 29640
rect 256516 27072 256568 27124
rect 400220 27072 400272 27124
rect 256424 27004 256476 27056
rect 407120 27004 407172 27056
rect 244740 26936 244792 26988
rect 447140 26936 447192 26988
rect 247592 26868 247644 26920
rect 471980 26868 472032 26920
rect 232320 25916 232372 25968
rect 280160 25916 280212 25968
rect 232228 25848 232280 25900
rect 284300 25848 284352 25900
rect 235080 25780 235132 25832
rect 311900 25780 311952 25832
rect 234988 25712 235040 25764
rect 318800 25712 318852 25764
rect 240600 25644 240652 25696
rect 390560 25644 390612 25696
rect 243360 25576 243412 25628
rect 425060 25576 425112 25628
rect 254400 25508 254452 25560
rect 567200 25508 567252 25560
rect 246120 24420 246172 24472
rect 463700 24420 463752 24472
rect 247316 24352 247368 24404
rect 473360 24352 473412 24404
rect 247408 24284 247460 24336
rect 477500 24284 477552 24336
rect 247500 24216 247552 24268
rect 481640 24216 481692 24268
rect 248972 24148 249024 24200
rect 490012 24148 490064 24200
rect 248880 24080 248932 24132
rect 496820 24080 496872 24132
rect 244924 23060 244976 23112
rect 386420 23060 386472 23112
rect 241704 22992 241756 23044
rect 407212 22992 407264 23044
rect 244556 22924 244608 22976
rect 441620 22924 441672 22976
rect 244648 22856 244700 22908
rect 448520 22856 448572 22908
rect 245936 22788 245988 22840
rect 456892 22788 456944 22840
rect 246028 22720 246080 22772
rect 459560 22720 459612 22772
rect 236460 21700 236512 21752
rect 335360 21700 335412 21752
rect 236368 21632 236420 21684
rect 339500 21632 339552 21684
rect 237932 21564 237984 21616
rect 349160 21564 349212 21616
rect 237840 21496 237892 21548
rect 357532 21496 357584 21548
rect 239220 21428 239272 21480
rect 371240 21428 371292 21480
rect 239128 21360 239180 21412
rect 374000 21360 374052 21412
rect 3424 20612 3476 20664
rect 199384 20612 199436 20664
rect 232136 20204 232188 20256
rect 285680 20204 285732 20256
rect 233608 20136 233660 20188
rect 296720 20136 296772 20188
rect 234896 20068 234948 20120
rect 314660 20068 314712 20120
rect 236276 20000 236328 20052
rect 332692 20000 332744 20052
rect 255412 19932 255464 19984
rect 578240 19932 578292 19984
rect 230848 19116 230900 19168
rect 267832 19116 267884 19168
rect 233884 19048 233936 19100
rect 271880 19048 271932 19100
rect 232044 18980 232096 19032
rect 278780 18980 278832 19032
rect 231952 18912 232004 18964
rect 282920 18912 282972 18964
rect 233516 18844 233568 18896
rect 303620 18844 303672 18896
rect 240508 18776 240560 18828
rect 396080 18776 396132 18828
rect 243268 18708 243320 18760
rect 418160 18708 418212 18760
rect 254216 18640 254268 18692
rect 563060 18640 563112 18692
rect 254308 18572 254360 18624
rect 569960 18572 570012 18624
rect 240416 17552 240468 17604
rect 397460 17552 397512 17604
rect 251548 17484 251600 17536
rect 527180 17484 527232 17536
rect 251640 17416 251692 17468
rect 534080 17416 534132 17468
rect 253020 17348 253072 17400
rect 545120 17348 545172 17400
rect 252836 17280 252888 17332
rect 547880 17280 547932 17332
rect 252928 17212 252980 17264
rect 552020 17212 552072 17264
rect 239036 16260 239088 16312
rect 376024 16260 376076 16312
rect 248604 16192 248656 16244
rect 495440 16192 495492 16244
rect 198740 16124 198792 16176
rect 225328 16124 225380 16176
rect 248696 16124 248748 16176
rect 498936 16124 498988 16176
rect 123024 16056 123076 16108
rect 219900 16056 219952 16108
rect 248788 16056 248840 16108
rect 502984 16056 503036 16108
rect 114008 15988 114060 16040
rect 218428 15988 218480 16040
rect 249892 15988 249944 16040
rect 509608 15988 509660 16040
rect 85672 15920 85724 15972
rect 210516 15920 210568 15972
rect 250076 15920 250128 15972
rect 513380 15920 513432 15972
rect 60832 15852 60884 15904
rect 211896 15852 211948 15904
rect 249984 15852 250036 15904
rect 517152 15852 517204 15904
rect 56784 14832 56836 14884
rect 214472 14832 214524 14884
rect 45008 14764 45060 14816
rect 212816 14764 212868 14816
rect 238944 14764 238996 14816
rect 369400 14764 369452 14816
rect 41880 14696 41932 14748
rect 211160 14696 211212 14748
rect 246948 14696 247000 14748
rect 462320 14696 462372 14748
rect 38384 14628 38436 14680
rect 212908 14628 212960 14680
rect 245844 14628 245896 14680
rect 465816 14628 465868 14680
rect 34520 14560 34572 14612
rect 211804 14560 211856 14612
rect 247040 14560 247092 14612
rect 473452 14560 473504 14612
rect 22560 14492 22612 14544
rect 211344 14492 211396 14544
rect 247224 14492 247276 14544
rect 476488 14492 476540 14544
rect 17960 14424 18012 14476
rect 211436 14424 211488 14476
rect 247132 14424 247184 14476
rect 481732 14424 481784 14476
rect 133144 13540 133196 13592
rect 215668 13540 215720 13592
rect 73344 13472 73396 13524
rect 215760 13472 215812 13524
rect 69848 13404 69900 13456
rect 215852 13404 215904 13456
rect 237748 13404 237800 13456
rect 351184 13404 351236 13456
rect 59360 13336 59412 13388
rect 214196 13336 214248 13388
rect 243176 13336 243228 13388
rect 430856 13336 430908 13388
rect 56048 13268 56100 13320
rect 214380 13268 214432 13320
rect 244280 13268 244332 13320
rect 440332 13268 440384 13320
rect 52552 13200 52604 13252
rect 214288 13200 214340 13252
rect 244464 13200 244516 13252
rect 445024 13200 445076 13252
rect 8760 13132 8812 13184
rect 210240 13132 210292 13184
rect 244372 13132 244424 13184
rect 448612 13132 448664 13184
rect 3608 13064 3660 13116
rect 210148 13064 210200 13116
rect 245660 13064 245712 13116
rect 459192 13064 459244 13116
rect 230756 12180 230808 12232
rect 264980 12180 265032 12232
rect 114744 12112 114796 12164
rect 218336 12112 218388 12164
rect 236184 12112 236236 12164
rect 330392 12112 330444 12164
rect 111616 12044 111668 12096
rect 218244 12044 218296 12096
rect 257436 12044 257488 12096
rect 415400 12044 415452 12096
rect 15936 11976 15988 12028
rect 178684 11976 178736 12028
rect 178776 11976 178828 12028
rect 212632 11976 212684 12028
rect 241520 11976 241572 12028
rect 406016 11976 406068 12028
rect 36728 11908 36780 11960
rect 212724 11908 212776 11960
rect 241612 11908 241664 11960
rect 409144 11908 409196 11960
rect 33600 11840 33652 11892
rect 213368 11840 213420 11892
rect 242992 11840 243044 11892
rect 420184 11840 420236 11892
rect 26240 11772 26292 11824
rect 211528 11772 211580 11824
rect 243084 11772 243136 11824
rect 423772 11772 423824 11824
rect 21824 11704 21876 11756
rect 211252 11704 211304 11756
rect 220820 11704 220872 11756
rect 221372 11704 221424 11756
rect 242900 11704 242952 11756
rect 426808 11704 426860 11756
rect 186964 10752 187016 10804
rect 218980 10752 219032 10804
rect 159364 10684 159416 10736
rect 218796 10684 218848 10736
rect 97448 10616 97500 10668
rect 216864 10616 216916 10668
rect 237656 10616 237708 10668
rect 359464 10616 359516 10668
rect 93952 10548 94004 10600
rect 217232 10548 217284 10600
rect 238852 10548 238904 10600
rect 370136 10548 370188 10600
rect 89904 10480 89956 10532
rect 217508 10480 217560 10532
rect 238760 10480 238812 10532
rect 374092 10480 374144 10532
rect 79232 10412 79284 10464
rect 215484 10412 215536 10464
rect 241428 10412 241480 10464
rect 390652 10412 390704 10464
rect 75920 10344 75972 10396
rect 215576 10344 215628 10396
rect 240324 10344 240376 10396
rect 395344 10344 395396 10396
rect 11152 10276 11204 10328
rect 188344 10276 188396 10328
rect 252744 10276 252796 10328
rect 553768 10276 553820 10328
rect 125876 9392 125928 9444
rect 215392 9392 215444 9444
rect 69112 9324 69164 9376
rect 216220 9324 216272 9376
rect 62028 9256 62080 9308
rect 214748 9256 214800 9308
rect 234804 9256 234856 9308
rect 324412 9256 324464 9308
rect 58440 9188 58492 9240
rect 214012 9188 214064 9240
rect 236092 9188 236144 9240
rect 338672 9188 338724 9240
rect 54944 9120 54996 9172
rect 214104 9120 214156 9172
rect 236000 9120 236052 9172
rect 342168 9120 342220 9172
rect 7656 9052 7708 9104
rect 209964 9052 210016 9104
rect 237472 9052 237524 9104
rect 349252 9052 349304 9104
rect 2872 8984 2924 9036
rect 209872 8984 209924 9036
rect 237380 8984 237432 9036
rect 352840 8984 352892 9036
rect 1676 8916 1728 8968
rect 210056 8916 210108 8968
rect 237564 8916 237616 8968
rect 356336 8916 356388 8968
rect 158904 7896 158956 7948
rect 222660 7896 222712 7948
rect 233332 7896 233384 7948
rect 303160 7896 303212 7948
rect 155408 7828 155460 7880
rect 220084 7828 220136 7880
rect 233240 7828 233292 7880
rect 306748 7828 306800 7880
rect 151912 7760 151964 7812
rect 221004 7760 221056 7812
rect 234620 7760 234672 7812
rect 317328 7760 317380 7812
rect 148324 7692 148376 7744
rect 221188 7692 221240 7744
rect 235908 7692 235960 7744
rect 320916 7692 320968 7744
rect 144736 7624 144788 7676
rect 221096 7624 221148 7676
rect 248512 7624 248564 7676
rect 492312 7624 492364 7676
rect 141240 7556 141292 7608
rect 221280 7556 221332 7608
rect 251456 7556 251508 7608
rect 529020 7556 529072 7608
rect 197912 6468 197964 6520
rect 225144 6468 225196 6520
rect 231860 6468 231912 6520
rect 285404 6468 285456 6520
rect 187332 6400 187384 6452
rect 223948 6400 224000 6452
rect 240140 6400 240192 6452
rect 388260 6400 388312 6452
rect 183744 6332 183796 6384
rect 223856 6332 223908 6384
rect 256332 6332 256384 6384
rect 562048 6332 562100 6384
rect 180248 6264 180300 6316
rect 223764 6264 223816 6316
rect 254032 6264 254084 6316
rect 566832 6264 566884 6316
rect 128176 6196 128228 6248
rect 219808 6196 219860 6248
rect 253940 6196 253992 6248
rect 569132 6196 569184 6248
rect 6460 6128 6512 6180
rect 209044 6128 209096 6180
rect 254124 6128 254176 6180
rect 572720 6128 572772 6180
rect 201592 5380 201644 5432
rect 225512 5380 225564 5432
rect 176752 5312 176804 5364
rect 224408 5312 224460 5364
rect 169576 5244 169628 5296
rect 222568 5244 222620 5296
rect 166080 5176 166132 5228
rect 223488 5176 223540 5228
rect 230664 5176 230716 5228
rect 262956 5176 263008 5228
rect 162492 5108 162544 5160
rect 222384 5108 222436 5160
rect 249800 5108 249852 5160
rect 519544 5108 519596 5160
rect 157800 5040 157852 5092
rect 222476 5040 222528 5092
rect 251364 5040 251416 5092
rect 525432 5040 525484 5092
rect 150624 4972 150676 5024
rect 220912 4972 220964 5024
rect 251272 4972 251324 5024
rect 533712 4972 533764 5024
rect 143540 4904 143592 4956
rect 221648 4904 221700 4956
rect 251180 4904 251232 4956
rect 537208 4904 537260 4956
rect 126980 4836 127032 4888
rect 219716 4836 219768 4888
rect 229376 4836 229428 4888
rect 247592 4836 247644 4888
rect 252652 4836 252704 4888
rect 547880 4836 547932 4888
rect 19432 4768 19484 4820
rect 203524 4768 203576 4820
rect 205088 4768 205140 4820
rect 225788 4768 225840 4820
rect 229468 4768 229520 4820
rect 252376 4768 252428 4820
rect 252560 4768 252612 4820
rect 554964 4768 555016 4820
rect 230572 4156 230624 4208
rect 186136 4088 186188 4140
rect 224316 4088 224368 4140
rect 227904 4088 227956 4140
rect 229836 4088 229888 4140
rect 182548 4020 182600 4072
rect 209136 4020 209188 4072
rect 210976 4020 211028 4072
rect 227168 4020 227220 4072
rect 95148 3952 95200 4004
rect 141424 3952 141476 4004
rect 151820 3952 151872 4004
rect 153016 3952 153068 4004
rect 168380 3952 168432 4004
rect 207664 3952 207716 4004
rect 213368 3952 213420 4004
rect 226524 3952 226576 4004
rect 104532 3884 104584 3936
rect 159364 3884 159416 3936
rect 164884 3884 164936 3936
rect 213184 3884 213236 3936
rect 215668 3884 215720 3936
rect 225604 3884 225656 3936
rect 99840 3816 99892 3868
rect 155224 3816 155276 3868
rect 167184 3816 167236 3868
rect 215944 3816 215996 3868
rect 219256 3816 219308 3868
rect 222844 3816 222896 3868
rect 256240 4088 256292 4140
rect 259460 4088 259512 4140
rect 261760 3816 261812 3868
rect 276020 3816 276072 3868
rect 276756 3816 276808 3868
rect 299572 3816 299624 3868
rect 300768 3816 300820 3868
rect 418804 3816 418856 3868
rect 581000 3816 581052 3868
rect 77392 3748 77444 3800
rect 133144 3748 133196 3800
rect 136456 3748 136508 3800
rect 213276 3748 213328 3800
rect 214472 3748 214524 3800
rect 226892 3748 226944 3800
rect 256056 3748 256108 3800
rect 465172 3748 465224 3800
rect 108120 3680 108172 3732
rect 186964 3680 187016 3732
rect 196808 3680 196860 3732
rect 210424 3680 210476 3732
rect 212172 3680 212224 3732
rect 226616 3680 226668 3732
rect 228088 3680 228140 3732
rect 235816 3680 235868 3732
rect 257344 3680 257396 3732
rect 468668 3680 468720 3732
rect 132960 3612 133012 3664
rect 219624 3612 219676 3664
rect 227812 3612 227864 3664
rect 237012 3612 237064 3664
rect 237380 3612 237432 3664
rect 258264 3612 258316 3664
rect 258724 3612 258776 3664
rect 72608 3544 72660 3596
rect 125876 3544 125928 3596
rect 129372 3544 129424 3596
rect 219532 3544 219584 3596
rect 230112 3544 230164 3596
rect 244096 3544 244148 3596
rect 248420 3544 248472 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 44272 3476 44324 3528
rect 52460 3408 52512 3460
rect 53380 3408 53432 3460
rect 176660 3476 176712 3528
rect 177856 3476 177908 3528
rect 201500 3476 201552 3528
rect 202696 3476 202748 3528
rect 223948 3476 224000 3528
rect 226432 3476 226484 3528
rect 227536 3476 227588 3528
rect 227996 3476 228048 3528
rect 231124 3476 231176 3528
rect 232228 3476 232280 3528
rect 47860 3340 47912 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 20628 3272 20680 3324
rect 25504 3272 25556 3324
rect 178776 3408 178828 3460
rect 207756 3408 207808 3460
rect 229192 3408 229244 3460
rect 250444 3476 250496 3528
rect 251180 3476 251232 3528
rect 253480 3408 253532 3460
rect 256148 3544 256200 3596
rect 479340 3680 479392 3732
rect 480536 3612 480588 3664
rect 473360 3544 473412 3596
rect 474188 3544 474240 3596
rect 481640 3544 481692 3596
rect 482468 3544 482520 3596
rect 255964 3476 256016 3528
rect 491116 3476 491168 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 501788 3408 501840 3460
rect 229284 3340 229336 3392
rect 246396 3340 246448 3392
rect 249984 3340 250036 3392
rect 256700 3340 256752 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365812 3340 365864 3392
rect 367008 3340 367060 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 226340 3136 226392 3188
rect 228180 3136 228232 3188
rect 242164 3136 242216 3188
rect 245200 3136 245252 3188
rect 232504 3068 232556 3120
rect 238116 3068 238168 3120
rect 423680 960 423732 1012
rect 424968 960 425020 1012
rect 448520 960 448572 1012
rect 449808 960 449860 1012
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3344 565894 3372 566879
rect 3332 565888 3384 565894
rect 3332 565830 3384 565836
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553450 3188 553823
rect 3148 553444 3200 553450
rect 3148 553386 3200 553392
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3252 474774 3280 475623
rect 3240 474768 3292 474774
rect 3240 474710 3292 474716
rect 2870 462632 2926 462641
rect 2870 462567 2926 462576
rect 2884 462398 2912 462567
rect 2872 462392 2924 462398
rect 2872 462334 2924 462340
rect 3238 449576 3294 449585
rect 3238 449511 3294 449520
rect 3252 447846 3280 449511
rect 3436 447914 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 449886 3556 671191
rect 3606 658200 3662 658209
rect 3606 658135 3662 658144
rect 3516 449880 3568 449886
rect 3516 449822 3568 449828
rect 3620 448050 3648 658135
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3712 448118 3740 632023
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3700 448112 3752 448118
rect 3700 448054 3752 448060
rect 3608 448044 3660 448050
rect 3608 447986 3660 447992
rect 3804 447982 3832 619103
rect 3882 606112 3938 606121
rect 3882 606047 3938 606056
rect 3896 449206 3924 606047
rect 3974 580000 4030 580009
rect 3974 579935 4030 579944
rect 3884 449200 3936 449206
rect 3884 449142 3936 449148
rect 3988 448186 4016 579935
rect 4066 514856 4122 514865
rect 4066 514791 4122 514800
rect 4080 464438 4108 514791
rect 4068 464432 4120 464438
rect 4068 464374 4120 464380
rect 6932 457502 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 22744 553444 22796 553450
rect 22744 553386 22796 553392
rect 14464 527196 14516 527202
rect 14464 527138 14516 527144
rect 10324 501016 10376 501022
rect 10324 500958 10376 500964
rect 10336 469946 10364 500958
rect 10324 469940 10376 469946
rect 10324 469882 10376 469888
rect 14476 460290 14504 527138
rect 22756 468518 22784 553386
rect 22744 468512 22796 468518
rect 22744 468454 22796 468460
rect 14464 460284 14516 460290
rect 14464 460226 14516 460232
rect 6920 457496 6972 457502
rect 6920 457438 6972 457444
rect 23492 448526 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 32404 565888 32456 565894
rect 32404 565830 32456 565836
rect 32416 472734 32444 565830
rect 32404 472728 32456 472734
rect 32404 472670 32456 472676
rect 40052 458862 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40684 474768 40736 474774
rect 40684 474710 40736 474716
rect 40696 471306 40724 474710
rect 40684 471300 40736 471306
rect 40684 471242 40736 471248
rect 71792 461718 71820 702986
rect 89180 700330 89208 703520
rect 105464 700398 105492 703520
rect 137848 700466 137876 703520
rect 154132 700534 154160 703520
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 170324 699718 170352 703520
rect 182824 700528 182876 700534
rect 182824 700470 182876 700476
rect 178684 700460 178736 700466
rect 178684 700402 178736 700408
rect 174544 700392 174596 700398
rect 174544 700334 174596 700340
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171784 699712 171836 699718
rect 171784 699654 171836 699660
rect 78586 636440 78642 636449
rect 78586 636375 78642 636384
rect 78310 635352 78366 635361
rect 78310 635287 78366 635296
rect 78218 633720 78274 633729
rect 78218 633655 78274 633664
rect 77758 632632 77814 632641
rect 77758 632567 77814 632576
rect 77772 523569 77800 632567
rect 78126 631000 78182 631009
rect 78126 630935 78182 630944
rect 77850 629640 77906 629649
rect 77850 629575 77906 629584
rect 77758 523560 77814 523569
rect 77758 523495 77814 523504
rect 77772 489666 77800 523495
rect 77864 520305 77892 629575
rect 78034 628008 78090 628017
rect 78034 627943 78090 627952
rect 77942 608696 77998 608705
rect 77942 608631 77998 608640
rect 77850 520296 77906 520305
rect 77850 520231 77906 520240
rect 77760 489660 77812 489666
rect 77760 489602 77812 489608
rect 77864 489462 77892 520231
rect 77956 498681 77984 608631
rect 78048 599962 78076 627943
rect 78140 600030 78168 630935
rect 78128 600024 78180 600030
rect 78128 599966 78180 599972
rect 78036 599956 78088 599962
rect 78036 599898 78088 599904
rect 78232 599826 78260 633655
rect 78220 599820 78272 599826
rect 78220 599762 78272 599768
rect 78324 587178 78352 635287
rect 78402 610056 78458 610065
rect 78402 609991 78458 610000
rect 78416 599758 78444 609991
rect 78494 607744 78550 607753
rect 78494 607679 78550 607688
rect 78404 599752 78456 599758
rect 78404 599694 78456 599700
rect 78508 599690 78536 607679
rect 78600 599894 78628 636375
rect 78588 599888 78640 599894
rect 78588 599830 78640 599836
rect 78496 599684 78548 599690
rect 78496 599626 78548 599632
rect 102874 597544 102930 597553
rect 102874 597479 102930 597488
rect 106186 597544 106242 597553
rect 106186 597479 106242 597488
rect 92478 597408 92534 597417
rect 92478 597343 92534 597352
rect 99286 597408 99342 597417
rect 99286 597343 99342 597352
rect 102046 597408 102102 597417
rect 102046 597343 102102 597352
rect 92492 596358 92520 597343
rect 94042 597000 94098 597009
rect 94042 596935 94098 596944
rect 97906 597000 97962 597009
rect 97906 596935 97908 596944
rect 79876 596352 79928 596358
rect 79876 596294 79928 596300
rect 92480 596352 92532 596358
rect 92480 596294 92532 596300
rect 79784 596284 79836 596290
rect 79784 596226 79836 596232
rect 78312 587172 78364 587178
rect 78312 587114 78364 587120
rect 78324 526561 78352 587114
rect 78494 526688 78550 526697
rect 78494 526623 78550 526632
rect 78310 526552 78366 526561
rect 78310 526487 78366 526496
rect 78310 523696 78366 523705
rect 78310 523631 78366 523640
rect 78126 520976 78182 520985
rect 78126 520911 78182 520920
rect 78034 499896 78090 499905
rect 78034 499831 78090 499840
rect 77942 498672 77998 498681
rect 77942 498607 77998 498616
rect 77852 489456 77904 489462
rect 77852 489398 77904 489404
rect 77956 474094 77984 498607
rect 78048 489598 78076 499831
rect 78140 489734 78168 520911
rect 78324 489802 78352 523631
rect 78402 498400 78458 498409
rect 78402 498335 78458 498344
rect 78312 489796 78364 489802
rect 78312 489738 78364 489744
rect 78128 489728 78180 489734
rect 78128 489670 78180 489676
rect 78036 489592 78088 489598
rect 78036 489534 78088 489540
rect 78416 489530 78444 498335
rect 78508 489870 78536 526623
rect 78586 517984 78642 517993
rect 78586 517919 78642 517928
rect 78496 489864 78548 489870
rect 78496 489806 78548 489812
rect 78404 489524 78456 489530
rect 78404 489466 78456 489472
rect 78600 489394 78628 517919
rect 78588 489388 78640 489394
rect 78588 489330 78640 489336
rect 79796 488442 79824 596226
rect 79888 488510 79916 596294
rect 94056 596290 94084 596935
rect 97960 596935 97962 596944
rect 97908 596906 97960 596912
rect 99300 596902 99328 597343
rect 100666 597136 100722 597145
rect 100666 597071 100722 597080
rect 100680 597038 100708 597071
rect 100668 597032 100720 597038
rect 100668 596974 100720 596980
rect 99288 596896 99340 596902
rect 99288 596838 99340 596844
rect 102060 596834 102088 597343
rect 102888 597310 102916 597479
rect 102876 597304 102928 597310
rect 102876 597246 102928 597252
rect 103426 597272 103482 597281
rect 103426 597207 103482 597216
rect 106094 597272 106150 597281
rect 106094 597207 106096 597216
rect 103440 597174 103468 597207
rect 106148 597207 106150 597216
rect 106096 597178 106148 597184
rect 103428 597168 103480 597174
rect 103428 597110 103480 597116
rect 104806 597136 104862 597145
rect 104806 597071 104808 597080
rect 104860 597071 104862 597080
rect 104808 597042 104860 597048
rect 102048 596828 102100 596834
rect 102048 596770 102100 596776
rect 95238 596320 95294 596329
rect 94044 596284 94096 596290
rect 95238 596255 95294 596264
rect 94044 596226 94096 596232
rect 95252 596222 95280 596255
rect 79968 596216 80020 596222
rect 79968 596158 80020 596164
rect 95240 596216 95292 596222
rect 95240 596158 95292 596164
rect 79876 488504 79928 488510
rect 79876 488446 79928 488452
rect 79784 488436 79836 488442
rect 79784 488378 79836 488384
rect 79980 488374 80008 596158
rect 106200 580310 106228 597479
rect 131026 597000 131082 597009
rect 131026 596935 131082 596944
rect 126886 596728 126942 596737
rect 126886 596663 126942 596672
rect 126900 596358 126928 596663
rect 131040 596426 131068 596935
rect 136546 596592 136602 596601
rect 136546 596527 136602 596536
rect 140686 596592 140742 596601
rect 140686 596527 140688 596536
rect 136560 596494 136588 596527
rect 140740 596527 140742 596536
rect 140688 596498 140740 596504
rect 136548 596488 136600 596494
rect 136548 596430 136600 596436
rect 131028 596420 131080 596426
rect 131028 596362 131080 596368
rect 126888 596352 126940 596358
rect 115846 596320 115902 596329
rect 115846 596255 115902 596264
rect 121366 596320 121422 596329
rect 126888 596294 126940 596300
rect 121366 596255 121368 596264
rect 115860 596222 115888 596255
rect 121420 596255 121422 596264
rect 121368 596226 121420 596232
rect 115848 596216 115900 596222
rect 115848 596158 115900 596164
rect 106188 580304 106240 580310
rect 106188 580246 106240 580252
rect 92940 488504 92992 488510
rect 92938 488472 92940 488481
rect 92992 488472 92994 488481
rect 92938 488407 92994 488416
rect 94226 488472 94282 488481
rect 94226 488407 94228 488416
rect 94280 488407 94282 488416
rect 95330 488472 95386 488481
rect 95330 488407 95386 488416
rect 97814 488472 97870 488481
rect 97814 488407 97870 488416
rect 98918 488472 98974 488481
rect 98918 488407 98974 488416
rect 100022 488472 100078 488481
rect 100022 488407 100078 488416
rect 101126 488472 101182 488481
rect 101126 488407 101182 488416
rect 102414 488472 102470 488481
rect 102414 488407 102470 488416
rect 104806 488472 104862 488481
rect 104806 488407 104862 488416
rect 105726 488472 105782 488481
rect 105726 488407 105782 488416
rect 94228 488378 94280 488384
rect 95344 488374 95372 488407
rect 79968 488368 80020 488374
rect 79968 488310 80020 488316
rect 95332 488368 95384 488374
rect 95332 488310 95384 488316
rect 97828 487218 97856 488407
rect 98932 487286 98960 488407
rect 100036 487354 100064 488407
rect 101140 487830 101168 488407
rect 101128 487824 101180 487830
rect 101128 487766 101180 487772
rect 102428 487422 102456 488407
rect 103426 488064 103482 488073
rect 104820 488034 104848 488407
rect 103426 487999 103482 488008
rect 104808 488028 104860 488034
rect 103440 487966 103468 487999
rect 104808 487970 104860 487976
rect 103428 487960 103480 487966
rect 103428 487902 103480 487908
rect 105740 487898 105768 488407
rect 106002 488200 106058 488209
rect 106002 488135 106058 488144
rect 111706 488200 111762 488209
rect 111706 488135 111762 488144
rect 105728 487892 105780 487898
rect 105728 487834 105780 487840
rect 102416 487416 102468 487422
rect 102416 487358 102468 487364
rect 100024 487348 100076 487354
rect 100024 487290 100076 487296
rect 98920 487280 98972 487286
rect 98920 487222 98972 487228
rect 97816 487212 97868 487218
rect 97816 487154 97868 487160
rect 106016 482390 106044 488135
rect 106004 482384 106056 482390
rect 106004 482326 106056 482332
rect 77944 474088 77996 474094
rect 77944 474030 77996 474036
rect 71780 461712 71832 461718
rect 71780 461654 71832 461660
rect 40040 458856 40092 458862
rect 40040 458798 40092 458804
rect 111720 449274 111748 488135
rect 115846 487248 115902 487257
rect 115846 487183 115902 487192
rect 121366 487248 121422 487257
rect 121366 487183 121422 487192
rect 126886 487248 126942 487257
rect 126886 487183 126942 487192
rect 131026 487248 131082 487257
rect 131026 487183 131082 487192
rect 136546 487248 136602 487257
rect 136546 487183 136602 487192
rect 140686 487248 140742 487257
rect 140686 487183 140742 487192
rect 115860 449342 115888 487183
rect 121380 467158 121408 487183
rect 126900 479602 126928 487183
rect 126888 479596 126940 479602
rect 126888 479538 126940 479544
rect 121368 467152 121420 467158
rect 121368 467094 121420 467100
rect 131040 461786 131068 487183
rect 136560 465866 136588 487183
rect 136548 465860 136600 465866
rect 136548 465802 136600 465808
rect 131028 461780 131080 461786
rect 131028 461722 131080 461728
rect 140700 449410 140728 487183
rect 171796 451994 171824 699654
rect 173254 596864 173310 596873
rect 173254 596799 173310 596808
rect 172244 596556 172296 596562
rect 172244 596498 172296 596504
rect 171876 596420 171928 596426
rect 171876 596362 171928 596368
rect 171784 451988 171836 451994
rect 171784 451930 171836 451936
rect 171888 449478 171916 596362
rect 171968 596284 172020 596290
rect 171968 596226 172020 596232
rect 171980 458930 172008 596226
rect 172152 596216 172204 596222
rect 172152 596158 172204 596164
rect 172060 580304 172112 580310
rect 172060 580246 172112 580252
rect 171968 458924 172020 458930
rect 171968 458866 172020 458872
rect 171876 449472 171928 449478
rect 171876 449414 171928 449420
rect 140688 449404 140740 449410
rect 140688 449346 140740 449352
rect 115848 449336 115900 449342
rect 115848 449278 115900 449284
rect 111708 449268 111760 449274
rect 111708 449210 111760 449216
rect 23480 448520 23532 448526
rect 23480 448462 23532 448468
rect 3976 448180 4028 448186
rect 3976 448122 4028 448128
rect 3792 447976 3844 447982
rect 3792 447918 3844 447924
rect 3424 447908 3476 447914
rect 3424 447850 3476 447856
rect 3240 447840 3292 447846
rect 3240 447782 3292 447788
rect 4988 446752 5040 446758
rect 4988 446694 5040 446700
rect 4804 446684 4856 446690
rect 4804 446626 4856 446632
rect 3516 446616 3568 446622
rect 3516 446558 3568 446564
rect 3240 443692 3292 443698
rect 3240 443634 3292 443640
rect 3148 423632 3200 423638
rect 3146 423600 3148 423609
rect 3200 423600 3202 423609
rect 3146 423535 3202 423544
rect 3252 410553 3280 443634
rect 3332 443216 3384 443222
rect 3332 443158 3384 443164
rect 3238 410544 3294 410553
rect 3238 410479 3294 410488
rect 3344 397497 3372 443158
rect 3424 443012 3476 443018
rect 3424 442954 3476 442960
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 2780 306264 2832 306270
rect 2778 306232 2780 306241
rect 2832 306232 2834 306241
rect 2778 306167 2834 306176
rect 3148 267708 3200 267714
rect 3148 267650 3200 267656
rect 3160 267209 3188 267650
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3056 215280 3108 215286
rect 3056 215222 3108 215228
rect 3068 214985 3096 215222
rect 3054 214976 3110 214985
rect 3054 214911 3110 214920
rect 2780 202700 2832 202706
rect 2780 202642 2832 202648
rect 2792 201929 2820 202642
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 3056 164212 3108 164218
rect 3056 164154 3108 164160
rect 3068 162897 3096 164154
rect 3054 162888 3110 162897
rect 3054 162823 3110 162832
rect 2780 149932 2832 149938
rect 2780 149874 2832 149880
rect 2792 149841 2820 149874
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3436 32473 3464 442954
rect 3528 58585 3556 446558
rect 3608 446344 3660 446350
rect 3608 446286 3660 446292
rect 3620 84697 3648 446286
rect 3792 445188 3844 445194
rect 3792 445130 3844 445136
rect 3700 445052 3752 445058
rect 3700 444994 3752 445000
rect 3712 136785 3740 444994
rect 3804 188873 3832 445130
rect 3884 445120 3936 445126
rect 3884 445062 3936 445068
rect 3896 241097 3924 445062
rect 4068 443284 4120 443290
rect 4068 443226 4120 443232
rect 3976 443148 4028 443154
rect 3976 443090 4028 443096
rect 3988 293185 4016 443090
rect 4080 345409 4108 443226
rect 4160 394460 4212 394466
rect 4160 394402 4212 394408
rect 4066 345400 4122 345409
rect 4066 345335 4122 345344
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3882 241088 3938 241097
rect 3882 241023 3938 241032
rect 3790 188864 3846 188873
rect 3790 188799 3846 188808
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 3606 84688 3662 84697
rect 3606 84623 3662 84632
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 394402
rect 4816 97782 4844 446626
rect 4896 443080 4948 443086
rect 4896 443022 4948 443028
rect 4908 149938 4936 443022
rect 5000 202706 5028 446694
rect 172072 446418 172100 580246
rect 172164 478378 172192 596158
rect 172256 486606 172284 596498
rect 173164 596352 173216 596358
rect 173164 596294 173216 596300
rect 172244 486600 172296 486606
rect 172244 486542 172296 486548
rect 173176 481098 173204 596294
rect 173268 485110 173296 596799
rect 173348 596488 173400 596494
rect 173348 596430 173400 596436
rect 173360 489258 173388 596430
rect 173348 489252 173400 489258
rect 173348 489194 173400 489200
rect 173256 485104 173308 485110
rect 173256 485046 173308 485052
rect 173164 481092 173216 481098
rect 173164 481034 173216 481040
rect 172152 478372 172204 478378
rect 172152 478314 172204 478320
rect 174556 457570 174584 700334
rect 178696 467294 178724 700402
rect 178684 467288 178736 467294
rect 178684 467230 178736 467236
rect 174544 457564 174596 457570
rect 174544 457506 174596 457512
rect 182836 453490 182864 700470
rect 202800 700466 202828 703520
rect 188896 700460 188948 700466
rect 188896 700402 188948 700408
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 184204 700324 184256 700330
rect 184204 700266 184256 700272
rect 188804 700324 188856 700330
rect 188804 700266 188856 700272
rect 182824 453484 182876 453490
rect 182824 453426 182876 453432
rect 184216 448254 184244 700266
rect 187330 637120 187386 637129
rect 187330 637055 187386 637064
rect 186778 636032 186834 636041
rect 186778 635967 186834 635976
rect 186686 630320 186742 630329
rect 186686 630255 186742 630264
rect 186700 520305 186728 630255
rect 186792 587178 186820 635967
rect 186870 634400 186926 634409
rect 186870 634335 186926 634344
rect 186884 599826 186912 634335
rect 187238 631680 187294 631689
rect 187238 631615 187294 631624
rect 187146 628688 187202 628697
rect 187146 628623 187202 628632
rect 187054 610328 187110 610337
rect 187054 610263 187110 610272
rect 186962 608424 187018 608433
rect 186962 608359 187018 608368
rect 186872 599820 186924 599826
rect 186872 599762 186924 599768
rect 186780 587172 186832 587178
rect 186780 587114 186832 587120
rect 186792 526017 186820 587114
rect 186778 526008 186834 526017
rect 186778 525943 186834 525952
rect 186884 524385 186912 599762
rect 186976 599690 187004 608359
rect 187068 599758 187096 610263
rect 187160 599962 187188 628623
rect 187252 600030 187280 631615
rect 187240 600024 187292 600030
rect 187240 599966 187292 599972
rect 187148 599956 187200 599962
rect 187148 599898 187200 599904
rect 187056 599752 187108 599758
rect 187056 599694 187108 599700
rect 186964 599684 187016 599690
rect 186964 599626 187016 599632
rect 186870 524376 186926 524385
rect 186870 524311 186926 524320
rect 186686 520296 186742 520305
rect 186686 520231 186742 520240
rect 186700 518894 186728 520231
rect 186700 518866 186912 518894
rect 186778 517576 186834 517585
rect 186778 517511 186834 517520
rect 186792 489394 186820 517511
rect 186884 489462 186912 518866
rect 186976 498409 187004 599626
rect 187068 500313 187096 599694
rect 187160 518673 187188 599898
rect 187252 521665 187280 599966
rect 187344 599894 187372 637055
rect 187422 633312 187478 633321
rect 187422 633247 187478 633256
rect 187332 599888 187384 599894
rect 187332 599830 187384 599836
rect 187344 527105 187372 599830
rect 187330 527096 187386 527105
rect 187330 527031 187386 527040
rect 187344 525842 187372 527031
rect 187332 525836 187384 525842
rect 187332 525778 187384 525784
rect 187436 523297 187464 633247
rect 187606 608696 187662 608705
rect 187606 608631 187662 608640
rect 187514 524376 187570 524385
rect 187514 524311 187570 524320
rect 187422 523288 187478 523297
rect 187422 523223 187478 523232
rect 187238 521656 187294 521665
rect 187238 521591 187294 521600
rect 187146 518664 187202 518673
rect 187146 518599 187202 518608
rect 187160 517585 187188 518599
rect 187146 517576 187202 517585
rect 187146 517511 187202 517520
rect 187054 500304 187110 500313
rect 187054 500239 187110 500248
rect 186962 498400 187018 498409
rect 186962 498335 187018 498344
rect 186976 489530 187004 498335
rect 187068 489598 187096 500239
rect 187252 489914 187280 521591
rect 187436 509234 187464 523223
rect 187160 489886 187280 489914
rect 187344 509206 187464 509234
rect 187160 489734 187188 489886
rect 187148 489728 187200 489734
rect 187148 489670 187200 489676
rect 187056 489592 187108 489598
rect 187056 489534 187108 489540
rect 186964 489524 187016 489530
rect 186964 489466 187016 489472
rect 186872 489456 186924 489462
rect 186872 489398 186924 489404
rect 186780 489388 186832 489394
rect 186780 489330 186832 489336
rect 186792 480254 186820 489330
rect 186884 488714 186912 489398
rect 186872 488708 186924 488714
rect 186872 488650 186924 488656
rect 186976 488578 187004 489466
rect 187068 488646 187096 489534
rect 187056 488640 187108 488646
rect 187056 488582 187108 488588
rect 186964 488572 187016 488578
rect 186964 488514 187016 488520
rect 186792 480226 187096 480254
rect 187068 449750 187096 480226
rect 187160 450770 187188 489670
rect 187344 489666 187372 509206
rect 187528 489802 187556 524311
rect 187620 498681 187648 608631
rect 188620 596352 188672 596358
rect 188620 596294 188672 596300
rect 188528 596216 188580 596222
rect 188528 596158 188580 596164
rect 188434 526008 188490 526017
rect 188434 525943 188490 525952
rect 187700 525836 187752 525842
rect 187700 525778 187752 525784
rect 187606 498672 187662 498681
rect 187606 498607 187662 498616
rect 187712 489870 187740 525778
rect 187700 489864 187752 489870
rect 187700 489806 187752 489812
rect 187516 489796 187568 489802
rect 187516 489738 187568 489744
rect 187332 489660 187384 489666
rect 187332 489602 187384 489608
rect 187240 488572 187292 488578
rect 187240 488514 187292 488520
rect 187148 450764 187200 450770
rect 187148 450706 187200 450712
rect 187252 450566 187280 488514
rect 187344 450838 187372 489602
rect 187424 488640 187476 488646
rect 187424 488582 187476 488588
rect 187332 450832 187384 450838
rect 187332 450774 187384 450780
rect 187436 450634 187464 488582
rect 187528 450702 187556 489738
rect 187608 488708 187660 488714
rect 187608 488650 187660 488656
rect 187516 450696 187568 450702
rect 187516 450638 187568 450644
rect 187424 450628 187476 450634
rect 187424 450570 187476 450576
rect 187240 450560 187292 450566
rect 187240 450502 187292 450508
rect 187056 449744 187108 449750
rect 187056 449686 187108 449692
rect 187620 449682 187648 488650
rect 187712 486538 187740 489806
rect 187700 486532 187752 486538
rect 187700 486474 187752 486480
rect 188448 450906 188476 525943
rect 188540 488442 188568 596158
rect 188632 488510 188660 596294
rect 188712 596284 188764 596290
rect 188712 596226 188764 596232
rect 188620 488504 188672 488510
rect 188620 488446 188672 488452
rect 188528 488436 188580 488442
rect 188528 488378 188580 488384
rect 188632 488238 188660 488446
rect 188620 488232 188672 488238
rect 188620 488174 188672 488180
rect 188724 488170 188752 596226
rect 188712 488164 188764 488170
rect 188712 488106 188764 488112
rect 188816 488102 188844 700266
rect 188804 488096 188856 488102
rect 188804 488038 188856 488044
rect 188436 450900 188488 450906
rect 188436 450842 188488 450848
rect 187608 449676 187660 449682
rect 187608 449618 187660 449624
rect 184204 448248 184256 448254
rect 184204 448190 184256 448196
rect 188908 446486 188936 700402
rect 218992 700398 219020 703520
rect 188988 700392 189040 700398
rect 188988 700334 189040 700340
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 189000 446554 189028 700334
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 281540 700324 281592 700330
rect 281540 700266 281592 700272
rect 207110 597544 207166 597553
rect 207110 597479 207166 597488
rect 208398 597544 208454 597553
rect 208398 597479 208454 597488
rect 210054 597544 210110 597553
rect 210054 597479 210110 597488
rect 211158 597544 211214 597553
rect 211158 597479 211214 597488
rect 212446 597544 212502 597553
rect 212446 597479 212502 597488
rect 213826 597544 213882 597553
rect 213826 597479 213882 597488
rect 214838 597544 214894 597553
rect 214838 597479 214894 597488
rect 215298 597544 215354 597553
rect 215298 597479 215354 597488
rect 215942 597544 215998 597553
rect 215942 597479 215998 597488
rect 226246 597544 226302 597553
rect 226246 597479 226302 597488
rect 235906 597544 235962 597553
rect 235906 597479 235962 597488
rect 245566 597544 245622 597553
rect 245566 597479 245622 597488
rect 251086 597544 251142 597553
rect 251086 597479 251142 597488
rect 204350 597136 204406 597145
rect 204350 597071 204406 597080
rect 202878 596456 202934 596465
rect 202878 596391 202934 596400
rect 202892 596358 202920 596391
rect 202880 596352 202932 596358
rect 202880 596294 202932 596300
rect 204258 596320 204314 596329
rect 204364 596290 204392 597071
rect 207124 596970 207152 597479
rect 207112 596964 207164 596970
rect 207112 596906 207164 596912
rect 204258 596255 204314 596264
rect 204352 596284 204404 596290
rect 204272 596222 204300 596255
rect 204352 596226 204404 596232
rect 207124 596222 207152 596906
rect 208412 596902 208440 597479
rect 210068 597038 210096 597479
rect 210056 597032 210108 597038
rect 210056 596974 210108 596980
rect 211068 597032 211120 597038
rect 211068 596974 211120 596980
rect 208400 596896 208452 596902
rect 208400 596838 208452 596844
rect 208412 596426 208440 596838
rect 208400 596420 208452 596426
rect 208400 596362 208452 596368
rect 211080 596358 211108 596974
rect 211172 596562 211200 597479
rect 212460 597310 212488 597479
rect 212448 597304 212500 597310
rect 212448 597246 212500 597252
rect 212460 596902 212488 597246
rect 213840 597174 213868 597479
rect 213828 597168 213880 597174
rect 213828 597110 213880 597116
rect 212448 596896 212500 596902
rect 212448 596838 212500 596844
rect 211160 596556 211212 596562
rect 211160 596498 211212 596504
rect 213840 596494 213868 597110
rect 214852 597106 214880 597479
rect 214840 597100 214892 597106
rect 214840 597042 214892 597048
rect 214852 596834 214880 597042
rect 214840 596828 214892 596834
rect 214840 596770 214892 596776
rect 213828 596488 213880 596494
rect 213828 596430 213880 596436
rect 211068 596352 211120 596358
rect 211068 596294 211120 596300
rect 204260 596216 204312 596222
rect 204260 596158 204312 596164
rect 207112 596216 207164 596222
rect 207112 596158 207164 596164
rect 215312 580378 215340 597479
rect 215956 597242 215984 597479
rect 215944 597236 215996 597242
rect 215944 597178 215996 597184
rect 215956 596698 215984 597178
rect 215944 596692 215996 596698
rect 215944 596634 215996 596640
rect 219438 596320 219494 596329
rect 219438 596255 219494 596264
rect 190000 580372 190052 580378
rect 190000 580314 190052 580320
rect 215300 580372 215352 580378
rect 215300 580314 215352 580320
rect 189908 580304 189960 580310
rect 189908 580246 189960 580252
rect 189078 498672 189134 498681
rect 189078 498607 189134 498616
rect 189092 450974 189120 498607
rect 189080 450968 189132 450974
rect 189080 450910 189132 450916
rect 189920 449546 189948 580246
rect 190012 449614 190040 580314
rect 219452 580310 219480 596255
rect 226260 581670 226288 597479
rect 231766 597272 231822 597281
rect 231766 597207 231822 597216
rect 226248 581664 226300 581670
rect 226248 581606 226300 581612
rect 231780 580310 231808 597207
rect 235920 580378 235948 597479
rect 241426 596864 241482 596873
rect 241426 596799 241482 596808
rect 241440 580446 241468 596799
rect 245580 580514 245608 597479
rect 251100 580582 251128 597479
rect 280988 596760 281040 596766
rect 280988 596702 281040 596708
rect 281000 596222 281028 596702
rect 280988 596216 281040 596222
rect 280988 596158 281040 596164
rect 251088 580576 251140 580582
rect 251088 580518 251140 580524
rect 245568 580508 245620 580514
rect 245568 580450 245620 580456
rect 241428 580440 241480 580446
rect 241428 580382 241480 580388
rect 235908 580372 235960 580378
rect 235908 580314 235960 580320
rect 219440 580304 219492 580310
rect 219440 580246 219492 580252
rect 231768 580304 231820 580310
rect 231768 580246 231820 580252
rect 253572 489252 253624 489258
rect 253572 489194 253624 489200
rect 218060 489184 218112 489190
rect 218060 489126 218112 489132
rect 204442 488472 204498 488481
rect 204442 488407 204444 488416
rect 204496 488407 204498 488416
rect 214838 488472 214894 488481
rect 214838 488407 214894 488416
rect 204444 488378 204496 488384
rect 202880 488232 202932 488238
rect 202878 488200 202880 488209
rect 202932 488200 202934 488209
rect 202878 488135 202934 488144
rect 204456 487490 204484 488378
rect 211158 488336 211214 488345
rect 211158 488271 211214 488280
rect 213734 488336 213790 488345
rect 213734 488271 213790 488280
rect 204904 488164 204956 488170
rect 204904 488106 204956 488112
rect 204444 487484 204496 487490
rect 204444 487426 204496 487432
rect 204916 487257 204944 488106
rect 211172 487830 211200 488271
rect 213748 487966 213776 488271
rect 214852 488034 214880 488407
rect 215390 488336 215446 488345
rect 215390 488271 215446 488280
rect 214840 488028 214892 488034
rect 214840 487970 214892 487976
rect 213736 487960 213788 487966
rect 213736 487902 213788 487908
rect 211160 487824 211212 487830
rect 211160 487766 211212 487772
rect 212448 487824 212500 487830
rect 212448 487766 212500 487772
rect 211802 487520 211858 487529
rect 211802 487455 211858 487464
rect 211816 487422 211844 487455
rect 212460 487422 212488 487766
rect 211804 487416 211856 487422
rect 210422 487384 210478 487393
rect 211804 487358 211856 487364
rect 212448 487416 212500 487422
rect 212448 487358 212500 487364
rect 210422 487319 210424 487328
rect 209056 487286 209084 487317
rect 210476 487319 210478 487328
rect 210424 487290 210476 487296
rect 209044 487280 209096 487286
rect 203522 487248 203578 487257
rect 203522 487183 203578 487192
rect 204902 487248 204958 487257
rect 204902 487183 204958 487192
rect 207662 487248 207718 487257
rect 207662 487183 207664 487192
rect 203536 459542 203564 487183
rect 203524 459536 203576 459542
rect 203524 459478 203576 459484
rect 204916 449818 204944 487183
rect 207716 487183 207718 487192
rect 209042 487248 209044 487257
rect 209096 487248 209098 487257
rect 209042 487183 209098 487192
rect 207664 487154 207716 487160
rect 207676 470558 207704 487154
rect 207664 470552 207716 470558
rect 207664 470494 207716 470500
rect 209056 463690 209084 487183
rect 210436 476814 210464 487290
rect 210424 476808 210476 476814
rect 210424 476750 210476 476756
rect 211816 471986 211844 487358
rect 213748 487286 213776 487902
rect 214852 487354 214880 487970
rect 215404 487898 215432 488271
rect 215392 487892 215444 487898
rect 215392 487834 215444 487840
rect 214840 487348 214892 487354
rect 214840 487290 214892 487296
rect 213736 487280 213788 487286
rect 213736 487222 213788 487228
rect 215404 487218 215432 487834
rect 216586 487248 216642 487257
rect 215392 487212 215444 487218
rect 216586 487183 216642 487192
rect 215392 487154 215444 487160
rect 215300 480956 215352 480962
rect 215300 480898 215352 480904
rect 211804 471980 211856 471986
rect 211804 471922 211856 471928
rect 214012 470620 214064 470626
rect 214012 470562 214064 470568
rect 209044 463684 209096 463690
rect 209044 463626 209096 463632
rect 204904 449812 204956 449818
rect 204904 449754 204956 449760
rect 190000 449608 190052 449614
rect 190000 449550 190052 449556
rect 189908 449540 189960 449546
rect 189908 449482 189960 449488
rect 214024 447370 214052 470562
rect 214196 460216 214248 460222
rect 214196 460158 214248 460164
rect 214012 447364 214064 447370
rect 214012 447306 214064 447312
rect 214208 447302 214236 460158
rect 214288 455524 214340 455530
rect 214288 455466 214340 455472
rect 214196 447296 214248 447302
rect 214196 447238 214248 447244
rect 213368 447160 213420 447166
rect 213368 447102 213420 447108
rect 188988 446548 189040 446554
rect 188988 446490 189040 446496
rect 188896 446480 188948 446486
rect 188896 446422 188948 446428
rect 172060 446412 172112 446418
rect 172060 446354 172112 446360
rect 213182 446312 213238 446321
rect 209136 446276 209188 446282
rect 213182 446247 213238 446256
rect 209136 446218 209188 446224
rect 5172 446140 5224 446146
rect 5172 446082 5224 446088
rect 5080 446072 5132 446078
rect 5080 446014 5132 446020
rect 5092 306270 5120 446014
rect 5184 358494 5212 446082
rect 208400 445800 208452 445806
rect 208400 445742 208452 445748
rect 196624 445596 196676 445602
rect 196624 445538 196676 445544
rect 98644 444508 98696 444514
rect 98644 444450 98696 444456
rect 13084 444440 13136 444446
rect 13084 444382 13136 444388
rect 13096 423638 13124 444382
rect 13084 423632 13136 423638
rect 13084 423574 13136 423580
rect 24860 398132 24912 398138
rect 24860 398074 24912 398080
rect 11058 396672 11114 396681
rect 11058 396607 11114 396616
rect 5172 358488 5224 358494
rect 5172 358430 5224 358436
rect 5080 306264 5132 306270
rect 5080 306206 5132 306212
rect 4988 202700 5040 202706
rect 4988 202642 5040 202648
rect 9680 177336 9732 177342
rect 9680 177278 9732 177284
rect 4896 149932 4948 149938
rect 4896 149874 4948 149880
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 4172 16546 5304 16574
rect 3608 13116 3660 13122
rect 3608 13058 3660 13064
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 1676 8968 1728 8974
rect 570 8936 626 8945
rect 1676 8910 1728 8916
rect 570 8871 626 8880
rect 584 480 612 8871
rect 1688 480 1716 8910
rect 2884 480 2912 8978
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 13058
rect 5276 480 5304 16546
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6472 480 6500 6122
rect 7668 480 7696 9046
rect 8772 480 8800 13126
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 177278
rect 11072 3534 11100 396607
rect 23480 338768 23532 338774
rect 23480 338710 23532 338716
rect 13818 177304 13874 177313
rect 13818 177239 13874 177248
rect 13832 16574 13860 177239
rect 23492 16574 23520 338710
rect 24872 16574 24900 398074
rect 25502 398032 25558 398041
rect 25502 397967 25558 397976
rect 13832 16546 14320 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 13542 14512 13598 14521
rect 13542 14447 13598 14456
rect 11152 10328 11204 10334
rect 11152 10270 11204 10276
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 10270
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 14447
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 22560 14544 22612 14550
rect 22560 14486 22612 14492
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 15936 12028 15988 12034
rect 15936 11970 15988 11976
rect 15948 480 15976 11970
rect 17038 11656 17094 11665
rect 17038 11591 17094 11600
rect 17052 480 17080 11591
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 14418
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19444 480 19472 4762
rect 20628 3324 20680 3330
rect 20628 3266 20680 3272
rect 20640 480 20668 3266
rect 21836 480 21864 11698
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 14486
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3330 25544 397967
rect 64878 396808 64934 396817
rect 40040 396772 40092 396778
rect 64878 396743 64934 396752
rect 40040 396714 40092 396720
rect 30380 395412 30432 395418
rect 30380 395354 30432 395360
rect 27620 395344 27672 395350
rect 27620 395286 27672 395292
rect 27710 395312 27766 395321
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 11766
rect 27632 6914 27660 395286
rect 27710 395247 27766 395256
rect 27724 16574 27752 395247
rect 28998 392592 29054 392601
rect 28998 392527 29054 392536
rect 29012 16574 29040 392527
rect 30392 16574 30420 395354
rect 35900 354000 35952 354006
rect 35900 353942 35952 353948
rect 31760 169040 31812 169046
rect 31760 168982 31812 168988
rect 31772 16574 31800 168982
rect 35912 16574 35940 353942
rect 38660 180124 38712 180130
rect 38660 180066 38712 180072
rect 38672 16574 38700 180066
rect 40052 16574 40080 396714
rect 52460 395480 52512 395486
rect 45558 395448 45614 395457
rect 52460 395422 52512 395428
rect 45558 395383 45614 395392
rect 42800 354068 42852 354074
rect 42800 354010 42852 354016
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 34520 14612 34572 14618
rect 34520 14554 34572 14560
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 33612 480 33640 11834
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 14554
rect 36004 480 36032 16546
rect 38384 14680 38436 14686
rect 38384 14622 38436 14628
rect 36728 11960 36780 11966
rect 36728 11902 36780 11908
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 11902
rect 38396 480 38424 14622
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 14748 41932 14754
rect 41880 14690 41932 14696
rect 41892 480 41920 14690
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 354010
rect 45572 16574 45600 395383
rect 49698 177440 49754 177449
rect 49698 177375 49754 177384
rect 49712 16574 49740 177375
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 45008 14816 45060 14822
rect 45008 14758 45060 14764
rect 44272 3528 44324 3534
rect 44272 3470 44324 3476
rect 44284 480 44312 3470
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 14758
rect 46676 480 46704 16546
rect 48502 13016 48558 13025
rect 48502 12951 48558 12960
rect 47860 3392 47912 3398
rect 47860 3334 47912 3340
rect 47872 480 47900 3334
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 12951
rect 50172 480 50200 16546
rect 51354 9072 51410 9081
rect 51354 9007 51410 9016
rect 51368 480 51396 9007
rect 52472 3466 52500 395422
rect 62120 354136 62172 354142
rect 62120 354078 62172 354084
rect 62132 16574 62160 354078
rect 63498 177576 63554 177585
rect 63498 177511 63554 177520
rect 63512 16574 63540 177511
rect 64892 16574 64920 396743
rect 67638 395584 67694 395593
rect 67638 395519 67694 395528
rect 77300 395548 77352 395554
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 60832 15904 60884 15910
rect 60832 15846 60884 15852
rect 56784 14884 56836 14890
rect 56784 14826 56836 14832
rect 56048 13320 56100 13326
rect 56048 13262 56100 13268
rect 52552 13252 52604 13258
rect 52552 13194 52604 13200
rect 52460 3460 52512 3466
rect 52460 3402 52512 3408
rect 52564 480 52592 13194
rect 54944 9172 54996 9178
rect 54944 9114 54996 9120
rect 53380 3460 53432 3466
rect 53380 3402 53432 3408
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3402
rect 54956 480 54984 9114
rect 56060 480 56088 13262
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 14826
rect 59360 13388 59412 13394
rect 59360 13330 59412 13336
rect 58440 9240 58492 9246
rect 58440 9182 58492 9188
rect 58452 480 58480 9182
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13330
rect 60844 480 60872 15846
rect 62028 9308 62080 9314
rect 62028 9250 62080 9256
rect 62040 480 62068 9250
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66718 13152 66774 13161
rect 66718 13087 66774 13096
rect 66732 480 66760 13087
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 395519
rect 77300 395490 77352 395496
rect 70400 354204 70452 354210
rect 70400 354146 70452 354152
rect 70412 16574 70440 354146
rect 74540 351212 74592 351218
rect 74540 351154 74592 351160
rect 74552 16574 74580 351154
rect 77312 16574 77340 395490
rect 92480 394052 92532 394058
rect 92480 393994 92532 394000
rect 91100 354340 91152 354346
rect 91100 354282 91152 354288
rect 86960 354272 87012 354278
rect 86960 354214 87012 354220
rect 80060 177404 80112 177410
rect 80060 177346 80112 177352
rect 80072 16574 80100 177346
rect 86972 16574 87000 354214
rect 88340 352572 88392 352578
rect 88340 352514 88392 352520
rect 88352 16574 88380 352514
rect 91112 16574 91140 354282
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 77312 16546 78168 16574
rect 80072 16546 80928 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 91112 16546 91600 16574
rect 69848 13456 69900 13462
rect 69848 13398 69900 13404
rect 69112 9376 69164 9382
rect 69112 9318 69164 9324
rect 69124 480 69152 9318
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 13398
rect 71516 480 71544 16546
rect 73344 13524 73396 13530
rect 73344 13466 73396 13472
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 72620 480 72648 3538
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 13466
rect 75012 480 75040 16546
rect 75920 10396 75972 10402
rect 75920 10338 75972 10344
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 10338
rect 77392 3800 77444 3806
rect 77392 3742 77444 3748
rect 77404 480 77432 3742
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 79232 10464 79284 10470
rect 79232 10406 79284 10412
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 10406
rect 80900 480 80928 16546
rect 85672 15972 85724 15978
rect 85672 15914 85724 15920
rect 84198 15872 84254 15881
rect 84198 15807 84254 15816
rect 81622 14648 81678 14657
rect 81622 14583 81678 14592
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 14583
rect 83278 10296 83334 10305
rect 83278 10231 83334 10240
rect 83292 480 83320 10231
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 15807
rect 85684 480 85712 15914
rect 86406 10432 86462 10441
rect 86406 10367 86462 10376
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 10367
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 89904 10532 89956 10538
rect 89904 10474 89956 10480
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 10474
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 393994
rect 98656 372570 98684 444450
rect 178682 398304 178738 398313
rect 171140 398268 171192 398274
rect 178682 398239 178738 398248
rect 171140 398210 171192 398216
rect 125600 398200 125652 398206
rect 125600 398142 125652 398148
rect 106280 396840 106332 396846
rect 106280 396782 106332 396788
rect 98644 372564 98696 372570
rect 98644 372506 98696 372512
rect 104900 355360 104952 355366
rect 102138 355328 102194 355337
rect 104900 355302 104952 355308
rect 102138 355263 102194 355272
rect 98000 354408 98052 354414
rect 98000 354350 98052 354356
rect 95240 82136 95292 82142
rect 95240 82078 95292 82084
rect 95252 16574 95280 82078
rect 98012 16574 98040 354350
rect 95252 16546 95832 16574
rect 98012 16546 98224 16574
rect 93952 10600 94004 10606
rect 93952 10542 94004 10548
rect 93964 480 93992 10542
rect 95148 4004 95200 4010
rect 95148 3946 95200 3952
rect 95160 480 95188 3946
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 97448 10668 97500 10674
rect 97448 10610 97500 10616
rect 97460 480 97488 10610
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 100758 10568 100814 10577
rect 100758 10503 100814 10512
rect 99840 3868 99892 3874
rect 99840 3810 99892 3816
rect 99852 480 99880 3810
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 10503
rect 102152 6914 102180 355263
rect 102232 178696 102284 178702
rect 102232 178638 102284 178644
rect 102244 16574 102272 178638
rect 104912 16574 104940 355302
rect 106292 16574 106320 396782
rect 118698 395720 118754 395729
rect 118698 395655 118754 395664
rect 115940 395616 115992 395622
rect 115940 395558 115992 395564
rect 109040 392624 109092 392630
rect 109040 392566 109092 392572
rect 102244 16546 103376 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 104532 3936 104584 3942
rect 104532 3878 104584 3884
rect 104544 480 104572 3878
rect 105740 480 105768 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 3732 108172 3738
rect 108120 3674 108172 3680
rect 108132 480 108160 3674
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 392566
rect 110420 355428 110472 355434
rect 110420 355370 110472 355376
rect 110432 16574 110460 355370
rect 111800 177472 111852 177478
rect 111800 177414 111852 177420
rect 111812 16574 111840 177414
rect 115952 16574 115980 395558
rect 117320 86284 117372 86290
rect 117320 86226 117372 86232
rect 110432 16546 110552 16574
rect 111812 16546 112392 16574
rect 115952 16546 116440 16574
rect 110524 480 110552 16546
rect 111616 12096 111668 12102
rect 111616 12038 111668 12044
rect 111628 480 111656 12038
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 16040 114060 16046
rect 114008 15982 114060 15988
rect 114020 480 114048 15982
rect 114744 12164 114796 12170
rect 114744 12106 114796 12112
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 12106
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 86226
rect 118712 3398 118740 395655
rect 120078 177712 120134 177721
rect 120078 177647 120134 177656
rect 120092 16574 120120 177647
rect 124220 177540 124272 177546
rect 124220 177482 124272 177488
rect 124232 16574 124260 177482
rect 120092 16546 120672 16574
rect 124232 16546 124720 16574
rect 118790 11792 118846 11801
rect 118790 11727 118846 11736
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 11727
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 123024 16108 123076 16114
rect 123024 16050 123076 16056
rect 122286 11928 122342 11937
rect 122286 11863 122342 11872
rect 122300 480 122328 11863
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16050
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 398142
rect 160100 397112 160152 397118
rect 160100 397054 160152 397060
rect 144920 397044 144972 397050
rect 144920 396986 144972 396992
rect 135260 396976 135312 396982
rect 135260 396918 135312 396924
rect 131120 396908 131172 396914
rect 131120 396850 131172 396856
rect 129740 394120 129792 394126
rect 129740 394062 129792 394068
rect 129752 16574 129780 394062
rect 131132 16574 131160 396850
rect 133880 394188 133932 394194
rect 133880 394130 133932 394136
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 125876 9444 125928 9450
rect 125876 9386 125928 9392
rect 125888 3602 125916 9386
rect 128176 6248 128228 6254
rect 128176 6190 128228 6196
rect 126980 4888 127032 4894
rect 126980 4830 127032 4836
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 126992 480 127020 4830
rect 128188 480 128216 6190
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 129384 480 129412 3538
rect 130580 480 130608 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 133144 13592 133196 13598
rect 133144 13534 133196 13540
rect 133156 3806 133184 13534
rect 133144 3800 133196 3806
rect 133144 3742 133196 3748
rect 132960 3664 133012 3670
rect 132960 3606 133012 3612
rect 132972 480 133000 3606
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 394130
rect 135272 480 135300 396918
rect 141424 395684 141476 395690
rect 141424 395626 141476 395632
rect 139398 393952 139454 393961
rect 139398 393887 139454 393896
rect 139412 16574 139440 393887
rect 139412 16546 139624 16574
rect 138846 16008 138902 16017
rect 138846 15943 138902 15952
rect 137650 6216 137706 6225
rect 137650 6151 137706 6160
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 136468 480 136496 3742
rect 137664 480 137692 6151
rect 138860 480 138888 15943
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141240 7608 141292 7614
rect 141240 7550 141292 7556
rect 141252 480 141280 7550
rect 141436 4010 141464 395626
rect 142160 351280 142212 351286
rect 142160 351222 142212 351228
rect 141424 4004 141476 4010
rect 141424 3946 141476 3952
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 351222
rect 144932 16574 144960 396986
rect 151818 396944 151874 396953
rect 151818 396879 151874 396888
rect 149060 352640 149112 352646
rect 149060 352582 149112 352588
rect 146300 46232 146352 46238
rect 146300 46174 146352 46180
rect 146312 16574 146340 46174
rect 149072 16574 149100 352582
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 149072 16546 149560 16574
rect 144736 7676 144788 7682
rect 144736 7618 144788 7624
rect 143540 4956 143592 4962
rect 143540 4898 143592 4904
rect 143552 480 143580 4898
rect 144748 480 144776 7618
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 148324 7744 148376 7750
rect 148324 7686 148376 7692
rect 148336 480 148364 7686
rect 149532 480 149560 16546
rect 150624 5024 150676 5030
rect 150624 4966 150676 4972
rect 150636 480 150664 4966
rect 151832 4010 151860 396879
rect 153198 352608 153254 352617
rect 153198 352543 153254 352552
rect 153212 16574 153240 352543
rect 155960 177608 156012 177614
rect 155960 177550 156012 177556
rect 155972 16574 156000 177550
rect 153212 16546 153792 16574
rect 155972 16546 156184 16574
rect 151912 7812 151964 7818
rect 151912 7754 151964 7760
rect 151820 4004 151872 4010
rect 151820 3946 151872 3952
rect 151924 3482 151952 7754
rect 153016 4004 153068 4010
rect 153016 3946 153068 3952
rect 151832 3454 151952 3482
rect 151832 480 151860 3454
rect 153028 480 153056 3946
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155222 14784 155278 14793
rect 155222 14719 155278 14728
rect 155236 3874 155264 14719
rect 155408 7880 155460 7886
rect 155408 7822 155460 7828
rect 155224 3868 155276 3874
rect 155224 3810 155276 3816
rect 155420 480 155448 7822
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 159364 10736 159416 10742
rect 159364 10678 159416 10684
rect 158904 7948 158956 7954
rect 158904 7890 158956 7896
rect 157800 5092 157852 5098
rect 157800 5034 157852 5040
rect 157812 480 157840 5034
rect 158916 480 158944 7890
rect 159376 3942 159404 10678
rect 159364 3936 159416 3942
rect 159364 3878 159416 3884
rect 160112 480 160140 397054
rect 160192 392692 160244 392698
rect 160192 392634 160244 392640
rect 160204 16574 160232 392634
rect 162860 46300 162912 46306
rect 162860 46242 162912 46248
rect 162872 16574 162900 46242
rect 171152 16574 171180 398210
rect 178040 394256 178092 394262
rect 178040 394198 178092 394204
rect 176660 354476 176712 354482
rect 176660 354418 176712 354424
rect 175278 351112 175334 351121
rect 175278 351047 175334 351056
rect 175292 16574 175320 351047
rect 160204 16546 161336 16574
rect 162872 16546 163728 16574
rect 171152 16546 172008 16574
rect 175292 16546 175504 16574
rect 161308 480 161336 16546
rect 162492 5160 162544 5166
rect 162492 5102 162544 5108
rect 162504 480 162532 5102
rect 163700 480 163728 16546
rect 170770 7576 170826 7585
rect 170770 7511 170826 7520
rect 169576 5296 169628 5302
rect 169576 5238 169628 5244
rect 166080 5228 166132 5234
rect 166080 5170 166132 5176
rect 164884 3936 164936 3942
rect 164884 3878 164936 3884
rect 164896 480 164924 3878
rect 166092 480 166120 5170
rect 168380 4004 168432 4010
rect 168380 3946 168432 3952
rect 167184 3868 167236 3874
rect 167184 3810 167236 3816
rect 167196 480 167224 3810
rect 168392 480 168420 3946
rect 169588 480 169616 5238
rect 170784 480 170812 7511
rect 171980 480 172008 16546
rect 174266 7712 174322 7721
rect 174266 7647 174322 7656
rect 173162 6352 173218 6361
rect 173162 6287 173218 6296
rect 173176 480 173204 6287
rect 174280 480 174308 7647
rect 175476 480 175504 16546
rect 176672 3534 176700 354418
rect 178052 16574 178080 394198
rect 178052 16546 178632 16574
rect 176752 5364 176804 5370
rect 176752 5306 176804 5312
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 176764 2666 176792 5306
rect 177856 3528 177908 3534
rect 177856 3470 177908 3476
rect 176672 2638 176792 2666
rect 176672 480 176700 2638
rect 177868 480 177896 3470
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 12034 178724 398239
rect 188342 398168 188398 398177
rect 188342 398103 188398 398112
rect 187698 392728 187754 392737
rect 187698 392663 187754 392672
rect 184940 355496 184992 355502
rect 184940 355438 184992 355444
rect 180800 354544 180852 354550
rect 180800 354486 180852 354492
rect 180812 16574 180840 354486
rect 180812 16546 181024 16574
rect 178684 12028 178736 12034
rect 178684 11970 178736 11976
rect 178776 12028 178828 12034
rect 178776 11970 178828 11976
rect 178788 3466 178816 11970
rect 180248 6316 180300 6322
rect 180248 6258 180300 6264
rect 178776 3460 178828 3466
rect 178776 3402 178828 3408
rect 180260 480 180288 6258
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 183744 6384 183796 6390
rect 183744 6326 183796 6332
rect 182548 4072 182600 4078
rect 182548 4014 182600 4020
rect 182560 480 182588 4014
rect 183756 480 183784 6326
rect 184952 480 184980 355438
rect 186964 10804 187016 10810
rect 186964 10746 187016 10752
rect 186136 4140 186188 4146
rect 186136 4082 186188 4088
rect 186148 480 186176 4082
rect 186976 3738 187004 10746
rect 187712 6914 187740 392663
rect 188356 10334 188384 398103
rect 193220 397724 193272 397730
rect 193220 397666 193272 397672
rect 189080 394324 189132 394330
rect 189080 394266 189132 394272
rect 189092 16574 189120 394266
rect 189092 16546 189304 16574
rect 188344 10328 188396 10334
rect 188344 10270 188396 10276
rect 187712 6886 188568 6914
rect 187332 6452 187384 6458
rect 187332 6394 187384 6400
rect 186964 3732 187016 3738
rect 186964 3674 187016 3680
rect 187344 480 187372 6394
rect 188540 480 188568 6886
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 192022 7848 192078 7857
rect 192022 7783 192078 7792
rect 190826 6488 190882 6497
rect 190826 6423 190882 6432
rect 190840 480 190868 6423
rect 192036 480 192064 7783
rect 193232 480 193260 397666
rect 194600 397180 194652 397186
rect 194600 397122 194652 397128
rect 194612 16574 194640 397122
rect 196636 164218 196664 445538
rect 199660 445460 199712 445466
rect 199660 445402 199712 445408
rect 196716 445392 196768 445398
rect 196716 445334 196768 445340
rect 196728 267714 196756 445334
rect 199568 445256 199620 445262
rect 199568 445198 199620 445204
rect 199476 444916 199528 444922
rect 199476 444858 199528 444864
rect 199384 443488 199436 443494
rect 199384 443430 199436 443436
rect 196716 267708 196768 267714
rect 196716 267650 196768 267656
rect 196624 164212 196676 164218
rect 196624 164154 196676 164160
rect 199396 20670 199424 443430
rect 199488 111790 199516 444858
rect 199580 215286 199608 445198
rect 199672 320142 199700 445402
rect 208412 445194 208440 445742
rect 208400 445188 208452 445194
rect 208400 445130 208452 445136
rect 209148 443972 209176 446218
rect 212078 446176 212134 446185
rect 212078 446111 212134 446120
rect 210422 446040 210478 446049
rect 210422 445975 210478 445984
rect 210238 445088 210294 445097
rect 210238 445023 210294 445032
rect 209686 444952 209742 444961
rect 209686 444887 209742 444896
rect 209502 444408 209558 444417
rect 209502 444343 209558 444352
rect 209332 444060 209452 444088
rect 209332 443972 209360 444060
rect 209424 443601 209452 444060
rect 209516 443972 209544 444343
rect 209700 443972 209728 444887
rect 210054 444680 210110 444689
rect 210054 444615 210110 444624
rect 209884 444060 210004 444088
rect 209884 443972 209912 444060
rect 209976 444009 210004 444060
rect 209962 444000 210018 444009
rect 210068 443972 210096 444615
rect 210252 443972 210280 445023
rect 210436 443972 210464 445975
rect 211068 445868 211120 445874
rect 211068 445810 211120 445816
rect 210792 445324 210844 445330
rect 210792 445266 210844 445272
rect 210606 444544 210662 444553
rect 210606 444479 210662 444488
rect 210620 443972 210648 444479
rect 210804 443972 210832 445266
rect 211080 445126 211108 445810
rect 211068 445120 211120 445126
rect 211068 445062 211120 445068
rect 211344 444780 211396 444786
rect 211344 444722 211396 444728
rect 210976 444712 211028 444718
rect 210976 444654 211028 444660
rect 210988 443972 211016 444654
rect 211172 444060 211292 444088
rect 211172 443972 211200 444060
rect 209962 443935 210018 443944
rect 211264 443737 211292 444060
rect 211356 443972 211384 444722
rect 211710 444136 211766 444145
rect 211540 444060 211660 444088
rect 211710 444071 211766 444080
rect 211540 443972 211568 444060
rect 211632 443873 211660 444060
rect 211724 443972 211752 444071
rect 211908 444060 212028 444088
rect 211908 443972 211936 444060
rect 211618 443864 211674 443873
rect 211618 443799 211674 443808
rect 211250 443728 211306 443737
rect 211250 443663 211306 443672
rect 209410 443592 209466 443601
rect 209410 443527 209466 443536
rect 212000 443465 212028 444060
rect 212092 443972 212120 446111
rect 212448 444848 212500 444854
rect 212448 444790 212500 444796
rect 212262 444136 212318 444145
rect 212262 444071 212318 444080
rect 212276 443972 212304 444071
rect 212460 443972 212488 444790
rect 212814 444136 212870 444145
rect 212644 444060 212764 444088
rect 212814 444071 212870 444080
rect 213000 444100 213052 444106
rect 212644 443972 212672 444060
rect 212540 443624 212592 443630
rect 212540 443566 212592 443572
rect 212552 443494 212580 443566
rect 212540 443488 212592 443494
rect 211986 443456 212042 443465
rect 212736 443465 212764 444060
rect 212828 443972 212856 444071
rect 213000 444042 213052 444048
rect 213012 443972 213040 444042
rect 213196 443972 213224 446247
rect 213380 443972 213408 447102
rect 213828 445936 213880 445942
rect 213828 445878 213880 445884
rect 213552 445188 213604 445194
rect 213552 445130 213604 445136
rect 213564 443972 213592 445130
rect 213840 445058 213868 445878
rect 213828 445052 213880 445058
rect 213828 444994 213880 445000
rect 213920 444644 213972 444650
rect 213920 444586 213972 444592
rect 213736 444576 213788 444582
rect 213736 444518 213788 444524
rect 213748 443972 213776 444518
rect 213932 443972 213960 444586
rect 214300 443972 214328 455466
rect 214472 455456 214524 455462
rect 214472 455398 214524 455404
rect 214484 443972 214512 455398
rect 214656 453348 214708 453354
rect 214656 453290 214708 453296
rect 214668 443972 214696 453290
rect 214840 451308 214892 451314
rect 214840 451250 214892 451256
rect 214852 443972 214880 451250
rect 215312 447370 215340 480898
rect 215484 479528 215536 479534
rect 215484 479470 215536 479476
rect 215392 472660 215444 472666
rect 215392 472602 215444 472608
rect 215024 447364 215076 447370
rect 215024 447306 215076 447312
rect 215300 447364 215352 447370
rect 215300 447306 215352 447312
rect 215036 443972 215064 447306
rect 215208 447296 215260 447302
rect 215208 447238 215260 447244
rect 215220 443972 215248 447238
rect 215404 443972 215432 472602
rect 215496 460934 215524 479470
rect 215668 474020 215720 474026
rect 215668 473962 215720 473968
rect 215496 460906 215616 460934
rect 215588 443972 215616 460906
rect 215680 445126 215708 473962
rect 216600 472802 216628 487183
rect 216772 486464 216824 486470
rect 216772 486406 216824 486412
rect 216680 482316 216732 482322
rect 216680 482258 216732 482264
rect 216588 472796 216640 472802
rect 216588 472738 216640 472744
rect 215852 464364 215904 464370
rect 215852 464306 215904 464312
rect 215760 461644 215812 461650
rect 215760 461586 215812 461592
rect 215668 445120 215720 445126
rect 215668 445062 215720 445068
rect 215772 443972 215800 461586
rect 215864 447302 215892 464306
rect 215944 453416 215996 453422
rect 215944 453358 215996 453364
rect 215852 447296 215904 447302
rect 215852 447238 215904 447244
rect 215956 443972 215984 453358
rect 216128 447364 216180 447370
rect 216128 447306 216180 447312
rect 216140 443972 216168 447306
rect 216312 447296 216364 447302
rect 216312 447238 216364 447244
rect 216324 443972 216352 447238
rect 216588 446004 216640 446010
rect 216588 445946 216640 445952
rect 216496 445120 216548 445126
rect 216496 445062 216548 445068
rect 216508 443972 216536 445062
rect 214196 443828 214248 443834
rect 214196 443770 214248 443776
rect 214208 443680 214236 443770
rect 216600 443698 216628 445946
rect 216692 443972 216720 482258
rect 216784 447302 216812 486406
rect 216956 483676 217008 483682
rect 216956 483618 217008 483624
rect 216864 463004 216916 463010
rect 216864 462946 216916 462952
rect 216772 447296 216824 447302
rect 216772 447238 216824 447244
rect 216876 443972 216904 462946
rect 216968 447250 216996 483618
rect 217140 475380 217192 475386
rect 217140 475322 217192 475328
rect 217152 447370 217180 475322
rect 217324 469872 217376 469878
rect 217324 469814 217376 469820
rect 217336 460934 217364 469814
rect 217508 465792 217560 465798
rect 217508 465734 217560 465740
rect 217520 460934 217548 465734
rect 217336 460906 217456 460934
rect 217520 460906 218008 460934
rect 217324 451920 217376 451926
rect 217324 451862 217376 451868
rect 217140 447364 217192 447370
rect 217140 447306 217192 447312
rect 216968 447222 217272 447250
rect 217048 445120 217100 445126
rect 217048 445062 217100 445068
rect 217060 443972 217088 445062
rect 217244 443972 217272 447222
rect 217336 445126 217364 451862
rect 217324 445120 217376 445126
rect 217324 445062 217376 445068
rect 217428 443972 217456 460906
rect 217600 447364 217652 447370
rect 217600 447306 217652 447312
rect 217612 443972 217640 447306
rect 217784 447296 217836 447302
rect 217784 447238 217836 447244
rect 217796 443972 217824 447238
rect 217980 443972 218008 460906
rect 218072 447370 218100 489126
rect 220084 488096 220136 488102
rect 220084 488038 220136 488044
rect 219808 487960 219860 487966
rect 219808 487902 219860 487908
rect 218244 478168 218296 478174
rect 218244 478110 218296 478116
rect 218152 476876 218204 476882
rect 218152 476818 218204 476824
rect 218060 447364 218112 447370
rect 218060 447306 218112 447312
rect 218164 443972 218192 476818
rect 218256 445126 218284 478110
rect 219624 468648 219676 468654
rect 219624 468590 219676 468596
rect 218336 468580 218388 468586
rect 218336 468522 218388 468528
rect 218244 445120 218296 445126
rect 218244 445062 218296 445068
rect 218348 443972 218376 468522
rect 218428 467220 218480 467226
rect 218428 467162 218480 467168
rect 218440 460934 218468 467162
rect 218440 460906 218560 460934
rect 218532 443972 218560 460906
rect 218612 460352 218664 460358
rect 218612 460294 218664 460300
rect 218624 447302 218652 460294
rect 219072 454708 219124 454714
rect 219072 454650 219124 454656
rect 218888 447364 218940 447370
rect 218888 447306 218940 447312
rect 218612 447296 218664 447302
rect 218612 447238 218664 447244
rect 218704 445120 218756 445126
rect 218704 445062 218756 445068
rect 218716 443972 218744 445062
rect 218900 443972 218928 447306
rect 219084 443972 219112 454650
rect 219440 447432 219492 447438
rect 219440 447374 219492 447380
rect 219256 447296 219308 447302
rect 219256 447238 219308 447244
rect 219268 443972 219296 447238
rect 219452 443972 219480 447374
rect 219636 443972 219664 468590
rect 219716 463208 219768 463214
rect 219716 463150 219768 463156
rect 219728 452198 219756 463150
rect 219716 452192 219768 452198
rect 219716 452134 219768 452140
rect 219820 445482 219848 487902
rect 219900 461848 219952 461854
rect 219900 461790 219952 461796
rect 219912 447438 219940 461790
rect 220096 460934 220124 488038
rect 230572 488028 230624 488034
rect 230572 487970 230624 487976
rect 222844 487484 222896 487490
rect 222844 487426 222896 487432
rect 220726 487248 220782 487257
rect 220726 487183 220782 487192
rect 220740 464574 220768 487183
rect 221464 484424 221516 484430
rect 221464 484366 221516 484372
rect 221372 467288 221424 467294
rect 221372 467230 221424 467236
rect 220728 464568 220780 464574
rect 220728 464510 220780 464516
rect 220096 460906 220216 460934
rect 219992 452192 220044 452198
rect 219992 452134 220044 452140
rect 219900 447432 219952 447438
rect 219900 447374 219952 447380
rect 219820 445454 219940 445482
rect 219912 444374 219940 445454
rect 219820 444346 219940 444374
rect 219820 443972 219848 444346
rect 220004 443972 220032 452134
rect 220082 444000 220138 444009
rect 220188 443972 220216 460906
rect 221004 458856 221056 458862
rect 221004 458798 221056 458804
rect 220820 457496 220872 457502
rect 220820 457438 220872 457444
rect 220728 451988 220780 451994
rect 220728 451930 220780 451936
rect 220544 446548 220596 446554
rect 220544 446490 220596 446496
rect 220360 446480 220412 446486
rect 220360 446422 220412 446428
rect 220268 444100 220320 444106
rect 220268 444042 220320 444048
rect 220082 443935 220138 443944
rect 217508 443828 217560 443834
rect 217508 443770 217560 443776
rect 214116 443652 214236 443680
rect 216588 443692 216640 443698
rect 214116 443564 214144 443652
rect 216588 443634 216640 443640
rect 212540 443430 212592 443436
rect 212722 443456 212778 443465
rect 211986 443391 212042 443400
rect 212722 443391 212778 443400
rect 215850 443456 215906 443465
rect 215850 443391 215852 443400
rect 215904 443391 215906 443400
rect 216586 443456 216642 443465
rect 217520 443426 217548 443770
rect 220096 443465 220124 443935
rect 220280 443562 220308 444042
rect 220372 443972 220400 446422
rect 220556 443972 220584 446490
rect 220740 443972 220768 451930
rect 220832 447234 220860 457438
rect 221016 447370 221044 458798
rect 221280 457564 221332 457570
rect 221280 457506 221332 457512
rect 221096 453484 221148 453490
rect 221096 453426 221148 453432
rect 221004 447364 221056 447370
rect 221004 447306 221056 447312
rect 220912 447296 220964 447302
rect 220912 447238 220964 447244
rect 220820 447228 220872 447234
rect 220820 447170 220872 447176
rect 220924 443972 220952 447238
rect 221108 443972 221136 453426
rect 221292 443972 221320 457506
rect 221384 447302 221412 467230
rect 221476 451314 221504 484366
rect 221556 461712 221608 461718
rect 221556 461654 221608 461660
rect 221464 451308 221516 451314
rect 221464 451250 221516 451256
rect 221372 447296 221424 447302
rect 221568 447284 221596 461654
rect 222200 448520 222252 448526
rect 222200 448462 222252 448468
rect 221648 448248 221700 448254
rect 221648 448190 221700 448196
rect 221372 447238 221424 447244
rect 221476 447256 221596 447284
rect 221476 443972 221504 447256
rect 221660 446214 221688 448190
rect 221832 447364 221884 447370
rect 221832 447306 221884 447312
rect 221648 446208 221700 446214
rect 221648 446150 221700 446156
rect 221660 443972 221688 446150
rect 221844 443972 221872 447306
rect 222016 447228 222068 447234
rect 222016 447170 222068 447176
rect 222028 443972 222056 447170
rect 222212 443972 222240 448462
rect 222856 448390 222884 487426
rect 226984 487416 227036 487422
rect 226984 487358 227036 487364
rect 226246 487248 226302 487257
rect 226246 487183 226302 487192
rect 224316 472728 224368 472734
rect 224316 472670 224368 472676
rect 223764 468512 223816 468518
rect 223764 468454 223816 468460
rect 222936 457292 222988 457298
rect 222936 457234 222988 457240
rect 222948 448526 222976 457234
rect 223028 456952 223080 456958
rect 223028 456894 223080 456900
rect 223040 449886 223068 456894
rect 223776 451274 223804 468454
rect 224224 464432 224276 464438
rect 224224 464374 224276 464380
rect 224040 460284 224092 460290
rect 224040 460226 224092 460232
rect 223856 456816 223908 456822
rect 223856 456758 223908 456764
rect 223684 451246 223804 451274
rect 223028 449880 223080 449886
rect 223028 449822 223080 449828
rect 222936 448520 222988 448526
rect 222936 448462 222988 448468
rect 222844 448384 222896 448390
rect 222844 448326 222896 448332
rect 223040 448202 223068 449822
rect 223120 449200 223172 449206
rect 223120 449142 223172 449148
rect 222764 448174 223068 448202
rect 222568 448044 222620 448050
rect 222568 447986 222620 447992
rect 222384 447908 222436 447914
rect 222384 447850 222436 447856
rect 222396 443972 222424 447850
rect 222580 443972 222608 447986
rect 222764 443972 222792 448174
rect 222936 448112 222988 448118
rect 222936 448054 222988 448060
rect 222948 443972 222976 448054
rect 223132 443972 223160 449142
rect 223488 448180 223540 448186
rect 223488 448122 223540 448128
rect 223304 447976 223356 447982
rect 223304 447918 223356 447924
rect 223316 447234 223344 447918
rect 223304 447228 223356 447234
rect 223304 447170 223356 447176
rect 223316 443972 223344 447170
rect 223500 443972 223528 448122
rect 223684 443972 223712 451246
rect 223868 443972 223896 456758
rect 224052 443972 224080 460226
rect 224236 451274 224264 464374
rect 224328 456822 224356 472670
rect 224500 471300 224552 471306
rect 224500 471242 224552 471248
rect 224512 460934 224540 471242
rect 224684 469940 224736 469946
rect 224684 469882 224736 469888
rect 224512 460906 224632 460934
rect 224316 456816 224368 456822
rect 224316 456758 224368 456764
rect 224236 451246 224448 451274
rect 224420 448633 224448 451246
rect 224406 448624 224462 448633
rect 224406 448559 224462 448568
rect 224224 447296 224276 447302
rect 224224 447238 224276 447244
rect 224236 443972 224264 447238
rect 224420 443972 224448 448559
rect 224604 443972 224632 460906
rect 224696 447302 224724 469882
rect 225604 462392 225656 462398
rect 225604 462334 225656 462340
rect 224776 447840 224828 447846
rect 224776 447782 224828 447788
rect 224684 447296 224736 447302
rect 224684 447238 224736 447244
rect 224788 443972 224816 447782
rect 225616 446826 225644 462334
rect 225694 454064 225750 454073
rect 225694 453999 225750 454008
rect 224960 446820 225012 446826
rect 224960 446762 225012 446768
rect 225604 446820 225656 446826
rect 225604 446762 225656 446768
rect 224972 443972 225000 446762
rect 225512 446004 225564 446010
rect 225512 445946 225564 445952
rect 225524 445534 225552 445946
rect 225512 445528 225564 445534
rect 225512 445470 225564 445476
rect 225144 444440 225196 444446
rect 225144 444382 225196 444388
rect 225156 443972 225184 444382
rect 225524 443972 225552 445470
rect 225708 444514 225736 453999
rect 226260 447846 226288 487183
rect 226996 448254 227024 487358
rect 229744 487348 229796 487354
rect 229744 487290 229796 487296
rect 227352 457496 227404 457502
rect 227352 457438 227404 457444
rect 226984 448248 227036 448254
rect 226984 448190 227036 448196
rect 226248 447840 226300 447846
rect 226248 447782 226300 447788
rect 227166 446584 227222 446593
rect 227166 446519 227222 446528
rect 226064 446140 226116 446146
rect 226064 446082 226116 446088
rect 225696 444508 225748 444514
rect 225696 444450 225748 444456
rect 225708 443972 225736 444450
rect 226076 443972 226104 446082
rect 226616 446072 226668 446078
rect 226616 446014 226668 446020
rect 226246 445904 226302 445913
rect 226246 445839 226302 445848
rect 226260 445466 226288 445839
rect 226248 445460 226300 445466
rect 226248 445402 226300 445408
rect 226260 443972 226288 445402
rect 226628 443972 226656 446014
rect 226984 445868 227036 445874
rect 226984 445810 227036 445816
rect 226800 445392 226852 445398
rect 226800 445334 226852 445340
rect 226812 444990 226840 445334
rect 226800 444984 226852 444990
rect 226800 444926 226852 444932
rect 226812 443972 226840 444926
rect 226996 443972 227024 445810
rect 227180 443972 227208 446519
rect 227364 445262 227392 457438
rect 228456 457224 228508 457230
rect 228456 457166 228508 457172
rect 228364 457088 228416 457094
rect 228364 457030 228416 457036
rect 227720 446752 227772 446758
rect 227720 446694 227772 446700
rect 227536 445800 227588 445806
rect 227536 445742 227588 445748
rect 227352 445256 227404 445262
rect 227352 445198 227404 445204
rect 227364 443972 227392 445198
rect 227548 443972 227576 445742
rect 227732 443972 227760 446694
rect 228088 445936 228140 445942
rect 228088 445878 228140 445884
rect 227904 445732 227956 445738
rect 227904 445674 227956 445680
rect 227916 445602 227944 445674
rect 227904 445596 227956 445602
rect 227904 445538 227956 445544
rect 227916 443972 227944 445538
rect 228100 443972 228128 445878
rect 228376 445618 228404 457030
rect 228468 445738 228496 457166
rect 229756 449886 229784 487290
rect 229836 487280 229888 487286
rect 229836 487222 229888 487228
rect 229848 451246 229876 487222
rect 229928 474088 229980 474094
rect 229928 474030 229980 474036
rect 229836 451240 229888 451246
rect 229836 451182 229888 451188
rect 229744 449880 229796 449886
rect 229744 449822 229796 449828
rect 229940 447098 229968 474030
rect 230584 460934 230612 487970
rect 232504 487892 232556 487898
rect 232504 487834 232556 487840
rect 231766 487248 231822 487257
rect 231766 487183 231822 487192
rect 231492 464500 231544 464506
rect 231492 464442 231544 464448
rect 230756 463072 230808 463078
rect 230756 463014 230808 463020
rect 230768 460934 230796 463014
rect 231504 460934 231532 464442
rect 230584 460906 230704 460934
rect 230768 460906 231256 460934
rect 231504 460906 231624 460934
rect 230676 451058 230704 460906
rect 230676 451030 231072 451058
rect 230848 450968 230900 450974
rect 230848 450910 230900 450916
rect 230480 448656 230532 448662
rect 230480 448598 230532 448604
rect 230296 448588 230348 448594
rect 230296 448530 230348 448536
rect 230112 447568 230164 447574
rect 230112 447510 230164 447516
rect 229928 447092 229980 447098
rect 229928 447034 229980 447040
rect 229190 446856 229246 446865
rect 229190 446791 229246 446800
rect 229006 446720 229062 446729
rect 228824 446684 228876 446690
rect 229006 446655 229062 446664
rect 228824 446626 228876 446632
rect 228640 446344 228692 446350
rect 228640 446286 228692 446292
rect 228456 445732 228508 445738
rect 228456 445674 228508 445680
rect 228376 445590 228496 445618
rect 228468 444922 228496 445590
rect 228456 444916 228508 444922
rect 228456 444858 228508 444864
rect 228468 443972 228496 444858
rect 228652 443972 228680 446286
rect 228836 443972 228864 446626
rect 229020 443972 229048 446655
rect 229204 443972 229232 446791
rect 229376 446616 229428 446622
rect 229376 446558 229428 446564
rect 229388 443972 229416 446558
rect 229742 446448 229798 446457
rect 229742 446383 229798 446392
rect 229560 445120 229612 445126
rect 229560 445062 229612 445068
rect 229572 444088 229600 445062
rect 229480 444060 229600 444088
rect 220268 443556 220320 443562
rect 220268 443498 220320 443504
rect 220082 443456 220138 443465
rect 216586 443391 216588 443400
rect 215852 443362 215904 443368
rect 216640 443391 216642 443400
rect 217508 443420 217560 443426
rect 216588 443362 216640 443368
rect 229480 443426 229508 444060
rect 229572 443972 229600 444060
rect 229756 443972 229784 446383
rect 230124 443972 230152 447510
rect 230308 443972 230336 448530
rect 230386 446584 230442 446593
rect 230386 446519 230442 446528
rect 230400 446282 230428 446519
rect 230388 446276 230440 446282
rect 230388 446218 230440 446224
rect 230492 443972 230520 448598
rect 230664 447092 230716 447098
rect 230664 447034 230716 447040
rect 230676 443972 230704 447034
rect 230860 443972 230888 450910
rect 231044 443972 231072 451030
rect 231228 443972 231256 460906
rect 231596 459542 231624 460906
rect 231584 459536 231636 459542
rect 231584 459478 231636 459484
rect 231398 445088 231454 445097
rect 231398 445023 231454 445032
rect 231412 443972 231440 445023
rect 231596 443972 231624 459478
rect 231780 447982 231808 487183
rect 232134 454336 232190 454345
rect 232134 454271 232190 454280
rect 231952 448384 232004 448390
rect 231952 448326 232004 448332
rect 231768 447976 231820 447982
rect 231768 447918 231820 447924
rect 231768 447432 231820 447438
rect 231768 447374 231820 447380
rect 231780 443972 231808 447374
rect 231964 443972 231992 448326
rect 232148 443972 232176 454271
rect 232516 448390 232544 487834
rect 232596 487824 232648 487830
rect 232596 487766 232648 487772
rect 232608 449818 232636 487766
rect 235906 487248 235962 487257
rect 235906 487183 235962 487192
rect 241426 487248 241482 487257
rect 241426 487183 241482 487192
rect 244646 487248 244702 487257
rect 249982 487248 250038 487257
rect 244646 487183 244702 487192
rect 244924 487212 244976 487218
rect 235264 486532 235316 486538
rect 235264 486474 235316 486480
rect 234620 482384 234672 482390
rect 234620 482326 234672 482332
rect 232686 454200 232742 454209
rect 232686 454135 232742 454144
rect 232596 449812 232648 449818
rect 232596 449754 232648 449760
rect 232504 448384 232556 448390
rect 232504 448326 232556 448332
rect 232608 448066 232636 449754
rect 232332 448038 232636 448066
rect 232332 443972 232360 448038
rect 232700 447250 232728 454135
rect 234632 451994 234660 482326
rect 235276 477426 235304 486474
rect 235264 477420 235316 477426
rect 235264 477362 235316 477368
rect 235276 476134 235304 477362
rect 234804 476128 234856 476134
rect 234804 476070 234856 476076
rect 235264 476128 235316 476134
rect 235264 476070 235316 476076
rect 234816 460934 234844 476070
rect 235920 474706 235948 487183
rect 240784 485172 240836 485178
rect 240784 485114 240836 485120
rect 236092 481024 236144 481030
rect 236092 480966 236144 480972
rect 235908 474700 235960 474706
rect 235908 474642 235960 474648
rect 235540 472796 235592 472802
rect 235540 472738 235592 472744
rect 235552 460934 235580 472738
rect 236104 460934 236132 480966
rect 238116 479732 238168 479738
rect 238116 479674 238168 479680
rect 236276 475448 236328 475454
rect 236276 475390 236328 475396
rect 234816 460906 234936 460934
rect 235552 460906 235856 460934
rect 236104 460906 236224 460934
rect 234712 454844 234764 454850
rect 234712 454786 234764 454792
rect 234620 451988 234672 451994
rect 234620 451930 234672 451936
rect 233976 451308 234028 451314
rect 233976 451250 234028 451256
rect 233792 450832 233844 450838
rect 233792 450774 233844 450780
rect 233424 450764 233476 450770
rect 233424 450706 233476 450712
rect 232780 449744 232832 449750
rect 232780 449686 232832 449692
rect 232516 447222 232728 447250
rect 232516 443972 232544 447222
rect 232792 444374 232820 449686
rect 233056 449676 233108 449682
rect 233056 449618 233108 449624
rect 232872 445868 232924 445874
rect 232872 445810 232924 445816
rect 232700 444346 232820 444374
rect 232700 443972 232728 444346
rect 232884 443972 232912 445810
rect 233068 443972 233096 449618
rect 233436 448322 233464 450706
rect 233424 448316 233476 448322
rect 233424 448258 233476 448264
rect 233240 446480 233292 446486
rect 233240 446422 233292 446428
rect 233252 443972 233280 446422
rect 233436 443972 233464 448258
rect 233804 448186 233832 450774
rect 233792 448180 233844 448186
rect 233792 448122 233844 448128
rect 233804 443972 233832 448122
rect 233988 443972 234016 451250
rect 234252 450900 234304 450906
rect 234252 450842 234304 450848
rect 234068 450696 234120 450702
rect 234068 450638 234120 450644
rect 234080 449857 234108 450638
rect 234066 449848 234122 449857
rect 234122 449806 234200 449834
rect 234066 449783 234122 449792
rect 234172 443972 234200 449806
rect 234264 449721 234292 450842
rect 234250 449712 234306 449721
rect 234250 449647 234306 449656
rect 234526 449712 234582 449721
rect 234526 449647 234582 449656
rect 234344 446140 234396 446146
rect 234344 446082 234396 446088
rect 234356 443972 234384 446082
rect 234540 443972 234568 449647
rect 234724 443972 234752 454786
rect 234908 443972 234936 460906
rect 235080 456068 235132 456074
rect 235080 456010 235132 456016
rect 235092 443972 235120 456010
rect 235264 454776 235316 454782
rect 235264 454718 235316 454724
rect 235276 443972 235304 454718
rect 235632 451988 235684 451994
rect 235632 451930 235684 451936
rect 235448 447432 235500 447438
rect 235448 447374 235500 447380
rect 235460 443972 235488 447374
rect 235644 443972 235672 451930
rect 235828 443972 235856 460906
rect 236000 445800 236052 445806
rect 236000 445742 236052 445748
rect 236012 443972 236040 445742
rect 236196 443972 236224 460906
rect 236288 445262 236316 475390
rect 237932 474088 237984 474094
rect 237932 474030 237984 474036
rect 236644 472796 236696 472802
rect 236644 472738 236696 472744
rect 236656 470558 236684 472738
rect 237472 471300 237524 471306
rect 237472 471242 237524 471248
rect 236644 470552 236696 470558
rect 236644 470494 236696 470500
rect 236368 457156 236420 457162
rect 236368 457098 236420 457104
rect 236276 445256 236328 445262
rect 236276 445198 236328 445204
rect 236380 443972 236408 457098
rect 236656 447134 236684 470494
rect 237012 464568 237064 464574
rect 237012 464510 237064 464516
rect 237024 460934 237052 464510
rect 237024 460906 237144 460934
rect 236920 449268 236972 449274
rect 236920 449210 236972 449216
rect 236736 447908 236788 447914
rect 236736 447850 236788 447856
rect 236564 447106 236684 447134
rect 236564 443972 236592 447106
rect 236748 443972 236776 447850
rect 236932 443972 236960 449210
rect 237116 443972 237144 460906
rect 237288 445256 237340 445262
rect 237288 445198 237340 445204
rect 237300 443972 237328 445198
rect 237484 443972 237512 471242
rect 237564 463684 237616 463690
rect 237564 463626 237616 463632
rect 237576 453150 237604 463626
rect 237748 455592 237800 455598
rect 237748 455534 237800 455540
rect 237564 453144 237616 453150
rect 237564 453086 237616 453092
rect 237760 444374 237788 455534
rect 237840 453144 237892 453150
rect 237840 453086 237892 453092
rect 237668 444346 237788 444374
rect 237668 443972 237696 444346
rect 237852 443972 237880 453086
rect 237944 445262 237972 474030
rect 238024 472728 238076 472734
rect 238024 472670 238076 472676
rect 238036 445806 238064 472670
rect 238128 463690 238156 479674
rect 238852 479664 238904 479670
rect 238852 479606 238904 479612
rect 238760 468512 238812 468518
rect 238760 468454 238812 468460
rect 238116 463684 238168 463690
rect 238116 463626 238168 463632
rect 238116 449744 238168 449750
rect 238116 449686 238168 449692
rect 238128 448526 238156 449686
rect 238208 449336 238260 449342
rect 238208 449278 238260 449284
rect 238116 448520 238168 448526
rect 238116 448462 238168 448468
rect 238116 446548 238168 446554
rect 238116 446490 238168 446496
rect 238024 445800 238076 445806
rect 238024 445742 238076 445748
rect 237932 445256 237984 445262
rect 237932 445198 237984 445204
rect 238128 444938 238156 446490
rect 238036 444910 238156 444938
rect 238036 443972 238064 444910
rect 238220 443972 238248 449278
rect 238392 447840 238444 447846
rect 238392 447782 238444 447788
rect 238404 443972 238432 447782
rect 238576 445256 238628 445262
rect 238576 445198 238628 445204
rect 238588 443972 238616 445198
rect 238772 443972 238800 468454
rect 238864 445262 238892 479606
rect 239404 476808 239456 476814
rect 239404 476750 239456 476756
rect 239036 469940 239088 469946
rect 239036 469882 239088 469888
rect 239048 451994 239076 469882
rect 239416 460834 239444 476750
rect 239496 467152 239548 467158
rect 239496 467094 239548 467100
rect 239404 460828 239456 460834
rect 239404 460770 239456 460776
rect 239036 451988 239088 451994
rect 239036 451930 239088 451936
rect 239416 447134 239444 460770
rect 239140 447106 239444 447134
rect 238852 445256 238904 445262
rect 238852 445198 238904 445204
rect 239140 443972 239168 447106
rect 239508 443972 239536 467094
rect 240324 464432 240376 464438
rect 240324 464374 240376 464380
rect 240048 451988 240100 451994
rect 240048 451930 240100 451936
rect 239588 449676 239640 449682
rect 239588 449618 239640 449624
rect 239600 448458 239628 449618
rect 239588 448452 239640 448458
rect 239588 448394 239640 448400
rect 239680 447976 239732 447982
rect 239680 447918 239732 447924
rect 239692 443972 239720 447918
rect 239864 445256 239916 445262
rect 239864 445198 239916 445204
rect 239876 443972 239904 445198
rect 240060 443972 240088 451930
rect 240232 445800 240284 445806
rect 240232 445742 240284 445748
rect 240244 443972 240272 445742
rect 240336 445262 240364 464374
rect 240508 463140 240560 463146
rect 240508 463082 240560 463088
rect 240520 456142 240548 463082
rect 240796 456794 240824 485114
rect 240876 479596 240928 479602
rect 240876 479538 240928 479544
rect 240612 456766 240824 456794
rect 240508 456136 240560 456142
rect 240508 456078 240560 456084
rect 240612 450786 240640 456766
rect 240428 450758 240640 450786
rect 240428 448254 240456 450758
rect 240416 448248 240468 448254
rect 240416 448190 240468 448196
rect 240324 445256 240376 445262
rect 240324 445198 240376 445204
rect 240428 443972 240456 448190
rect 240600 447636 240652 447642
rect 240600 447578 240652 447584
rect 240612 443972 240640 447578
rect 240888 447134 240916 479538
rect 241440 474706 241468 487183
rect 243544 486668 243596 486674
rect 243544 486610 243596 486616
rect 242164 482452 242216 482458
rect 242164 482394 242216 482400
rect 241612 476808 241664 476814
rect 241612 476750 241664 476756
rect 240968 474700 241020 474706
rect 240968 474642 241020 474648
rect 241428 474700 241480 474706
rect 241428 474642 241480 474648
rect 240796 447106 240916 447134
rect 240796 443972 240824 447106
rect 240980 443972 241008 474642
rect 241152 456136 241204 456142
rect 241152 456078 241204 456084
rect 241164 443972 241192 456078
rect 241624 451994 241652 476750
rect 242176 471986 242204 482394
rect 242256 474700 242308 474706
rect 242256 474642 242308 474648
rect 241704 471980 241756 471986
rect 241704 471922 241756 471928
rect 242164 471980 242216 471986
rect 242164 471922 242216 471928
rect 241612 451988 241664 451994
rect 241612 451930 241664 451936
rect 241520 449200 241572 449206
rect 241520 449142 241572 449148
rect 241336 445256 241388 445262
rect 241336 445198 241388 445204
rect 241348 443972 241376 445198
rect 241532 443972 241560 449142
rect 241716 443972 241744 471922
rect 242072 461780 242124 461786
rect 242072 461722 242124 461728
rect 241796 461712 241848 461718
rect 241796 461654 241848 461660
rect 241808 445262 241836 461654
rect 241888 447568 241940 447574
rect 241888 447510 241940 447516
rect 241796 445256 241848 445262
rect 241796 445198 241848 445204
rect 241900 443972 241928 447510
rect 242084 443972 242112 461722
rect 242268 443972 242296 474642
rect 243360 465860 243412 465866
rect 243360 465802 243412 465808
rect 243084 465724 243136 465730
rect 243084 465666 243136 465672
rect 243096 451994 243124 465666
rect 243176 452532 243228 452538
rect 243176 452474 243228 452480
rect 242624 451988 242676 451994
rect 242624 451930 242676 451936
rect 243084 451988 243136 451994
rect 243084 451930 243136 451936
rect 242440 445256 242492 445262
rect 242440 445198 242492 445204
rect 242452 443972 242480 445198
rect 242636 443972 242664 451930
rect 242992 451240 243044 451246
rect 242992 451182 243044 451188
rect 243004 443972 243032 451182
rect 243188 443972 243216 452474
rect 243372 443972 243400 465802
rect 243556 451246 243584 486610
rect 244660 485858 244688 487183
rect 249982 487183 250038 487192
rect 244924 487154 244976 487160
rect 243636 485852 243688 485858
rect 243636 485794 243688 485800
rect 244648 485852 244700 485858
rect 244648 485794 244700 485800
rect 243544 451240 243596 451246
rect 243544 451182 243596 451188
rect 243648 447134 243676 485794
rect 244936 476066 244964 487154
rect 247224 485104 247276 485110
rect 247224 485046 247276 485052
rect 248420 485104 248472 485110
rect 248420 485046 248472 485052
rect 246396 482384 246448 482390
rect 246396 482326 246448 482332
rect 244372 476060 244424 476066
rect 244372 476002 244424 476008
rect 244924 476060 244976 476066
rect 244924 476002 244976 476008
rect 243912 451988 243964 451994
rect 243912 451930 243964 451936
rect 243556 447106 243676 447134
rect 243556 443972 243584 447106
rect 243728 447092 243780 447098
rect 243728 447034 243780 447040
rect 243740 443972 243768 447034
rect 243924 443972 243952 451930
rect 244280 448792 244332 448798
rect 244280 448734 244332 448740
rect 244096 448724 244148 448730
rect 244096 448666 244148 448672
rect 244108 443972 244136 448666
rect 244292 443972 244320 448734
rect 244384 447506 244412 476002
rect 244924 474156 244976 474162
rect 244924 474098 244976 474104
rect 244556 467152 244608 467158
rect 244556 467094 244608 467100
rect 244568 460934 244596 467094
rect 244568 460906 244872 460934
rect 244464 455728 244516 455734
rect 244464 455670 244516 455676
rect 244372 447500 244424 447506
rect 244372 447442 244424 447448
rect 244476 443972 244504 455670
rect 244648 449404 244700 449410
rect 244648 449346 244700 449352
rect 244660 443972 244688 449346
rect 244740 447704 244792 447710
rect 244740 447646 244792 447652
rect 244752 447134 244780 447646
rect 244844 447250 244872 460906
rect 244936 449886 244964 474098
rect 246304 458992 246356 458998
rect 246304 458934 246356 458940
rect 245844 452056 245896 452062
rect 245844 451998 245896 452004
rect 244924 449880 244976 449886
rect 244924 449822 244976 449828
rect 244936 448798 244964 449822
rect 244924 448792 244976 448798
rect 244924 448734 244976 448740
rect 245752 447840 245804 447846
rect 245752 447782 245804 447788
rect 245568 447500 245620 447506
rect 245568 447442 245620 447448
rect 244844 447222 245240 447250
rect 244752 447106 244872 447134
rect 244844 443972 244872 447106
rect 245016 445868 245068 445874
rect 245016 445810 245068 445816
rect 245028 443972 245056 445810
rect 245212 443972 245240 447222
rect 245384 445936 245436 445942
rect 245384 445878 245436 445884
rect 245396 443972 245424 445878
rect 245580 443972 245608 447442
rect 245764 443972 245792 447782
rect 245856 447506 245884 451998
rect 246120 449608 246172 449614
rect 246120 449550 246172 449556
rect 245844 447500 245896 447506
rect 245844 447442 245896 447448
rect 245936 446412 245988 446418
rect 245936 446354 245988 446360
rect 245948 443972 245976 446354
rect 246132 443972 246160 449550
rect 246212 447772 246264 447778
rect 246212 447714 246264 447720
rect 246224 447098 246252 447714
rect 246316 447574 246344 458934
rect 246304 447568 246356 447574
rect 246304 447510 246356 447516
rect 246408 447386 246436 482326
rect 246488 478304 246540 478310
rect 246488 478246 246540 478252
rect 246500 447778 246528 478246
rect 246764 478236 246816 478242
rect 246764 478178 246816 478184
rect 246776 451274 246804 478178
rect 247040 458856 247092 458862
rect 247040 458798 247092 458804
rect 247052 452538 247080 458798
rect 247132 457020 247184 457026
rect 247132 456962 247184 456968
rect 247040 452532 247092 452538
rect 247040 452474 247092 452480
rect 246592 451246 246804 451274
rect 246488 447772 246540 447778
rect 246488 447714 246540 447720
rect 246316 447358 246436 447386
rect 246212 447092 246264 447098
rect 246212 447034 246264 447040
rect 246316 445874 246344 447358
rect 246592 447250 246620 451246
rect 246672 449268 246724 449274
rect 246672 449210 246724 449216
rect 246500 447222 246620 447250
rect 246396 446684 246448 446690
rect 246396 446626 246448 446632
rect 246304 445868 246356 445874
rect 246304 445810 246356 445816
rect 246408 444938 246436 446626
rect 246316 444910 246436 444938
rect 246316 443972 246344 444910
rect 246500 443972 246528 447222
rect 246684 443972 246712 449210
rect 247040 448792 247092 448798
rect 247040 448734 247092 448740
rect 246856 447500 246908 447506
rect 246856 447442 246908 447448
rect 246868 443972 246896 447442
rect 246948 446208 247000 446214
rect 246948 446150 247000 446156
rect 246960 445058 246988 446150
rect 246948 445052 247000 445058
rect 246948 444994 247000 445000
rect 247052 443972 247080 448734
rect 247144 445262 247172 456962
rect 247132 445256 247184 445262
rect 247132 445198 247184 445204
rect 247236 443972 247264 485046
rect 248144 452192 248196 452198
rect 248144 452134 248196 452140
rect 247408 451988 247460 451994
rect 247408 451930 247460 451936
rect 247316 449540 247368 449546
rect 247316 449482 247368 449488
rect 247328 447134 247356 449482
rect 247420 447250 247448 451930
rect 247420 447222 248000 447250
rect 247328 447106 247448 447134
rect 247420 443972 247448 447106
rect 247776 446956 247828 446962
rect 247776 446898 247828 446904
rect 247592 446616 247644 446622
rect 247592 446558 247644 446564
rect 247604 443972 247632 446558
rect 247788 443972 247816 446898
rect 247972 443972 248000 447222
rect 248156 443972 248184 452134
rect 248432 445262 248460 485046
rect 248512 478372 248564 478378
rect 248512 478314 248564 478320
rect 248328 445256 248380 445262
rect 248328 445198 248380 445204
rect 248420 445256 248472 445262
rect 248420 445198 248472 445204
rect 248340 443972 248368 445198
rect 248524 443972 248552 478314
rect 249800 458924 249852 458930
rect 249800 458866 249852 458872
rect 248696 454912 248748 454918
rect 248696 454854 248748 454860
rect 248708 449290 248736 454854
rect 249432 452124 249484 452130
rect 249432 452066 249484 452072
rect 248708 449262 249288 449290
rect 248696 449132 248748 449138
rect 248696 449074 248748 449080
rect 248708 443972 248736 449074
rect 248972 446820 249024 446826
rect 248972 446762 249024 446768
rect 248880 446208 248932 446214
rect 248880 446150 248932 446156
rect 248892 443972 248920 446150
rect 248984 443698 249012 446762
rect 249064 445256 249116 445262
rect 249064 445198 249116 445204
rect 249076 443972 249104 445198
rect 249260 443972 249288 449262
rect 249444 443972 249472 452066
rect 249616 448860 249668 448866
rect 249616 448802 249668 448808
rect 249628 443972 249656 448802
rect 249812 443972 249840 458866
rect 249892 449336 249944 449342
rect 249892 449278 249944 449284
rect 249904 447134 249932 449278
rect 249996 447710 250024 487183
rect 251640 483744 251692 483750
rect 251640 483686 251692 483692
rect 250996 481092 251048 481098
rect 250996 481034 251048 481040
rect 251008 460934 251036 481034
rect 251008 460906 251128 460934
rect 250168 455796 250220 455802
rect 250168 455738 250220 455744
rect 249984 447704 250036 447710
rect 249984 447646 250036 447652
rect 250180 447250 250208 455738
rect 250720 452328 250772 452334
rect 250720 452270 250772 452276
rect 250180 447222 250576 447250
rect 249904 447106 250024 447134
rect 249892 446004 249944 446010
rect 249892 445946 249944 445952
rect 249904 443766 249932 445946
rect 249996 443972 250024 447106
rect 250352 447024 250404 447030
rect 250352 446966 250404 446972
rect 250168 446888 250220 446894
rect 250168 446830 250220 446836
rect 250180 443972 250208 446830
rect 250364 443972 250392 446966
rect 250548 443972 250576 447222
rect 250732 443972 250760 452270
rect 250902 444136 250958 444145
rect 250902 444071 250958 444080
rect 250916 443972 250944 444071
rect 251100 443972 251128 460906
rect 251364 455864 251416 455870
rect 251364 455806 251416 455812
rect 251272 449404 251324 449410
rect 251272 449346 251324 449352
rect 251284 443972 251312 449346
rect 251376 447574 251404 455806
rect 251548 452260 251600 452266
rect 251548 452202 251600 452208
rect 251364 447568 251416 447574
rect 251364 447510 251416 447516
rect 251456 446820 251508 446826
rect 251456 446762 251508 446768
rect 251468 443972 251496 446762
rect 251560 444242 251588 452202
rect 251548 444236 251600 444242
rect 251548 444178 251600 444184
rect 251652 443972 251680 483686
rect 253584 460934 253612 489194
rect 254860 486600 254912 486606
rect 254860 486542 254912 486548
rect 253940 486532 253992 486538
rect 253940 486474 253992 486480
rect 253952 460934 253980 486474
rect 254872 460934 254900 486542
rect 253584 460906 253704 460934
rect 253952 460906 254072 460934
rect 254872 460906 254992 460934
rect 253296 458924 253348 458930
rect 253296 458866 253348 458872
rect 252652 456000 252704 456006
rect 252652 455942 252704 455948
rect 251732 455932 251784 455938
rect 251732 455874 251784 455880
rect 251744 446486 251772 455874
rect 252560 449540 252612 449546
rect 252560 449482 252612 449488
rect 252376 449472 252428 449478
rect 252376 449414 252428 449420
rect 252192 448928 252244 448934
rect 252192 448870 252244 448876
rect 251824 447568 251876 447574
rect 251824 447510 251876 447516
rect 251732 446480 251784 446486
rect 251732 446422 251784 446428
rect 251836 443972 251864 447510
rect 252008 444236 252060 444242
rect 252008 444178 252060 444184
rect 252020 443972 252048 444178
rect 252204 443972 252232 448870
rect 252388 443972 252416 449414
rect 252572 443972 252600 449482
rect 252664 447250 252692 455942
rect 253204 452396 253256 452402
rect 253204 452338 253256 452344
rect 252744 449336 252796 449342
rect 252744 449278 252796 449284
rect 252756 449138 252784 449278
rect 252744 449132 252796 449138
rect 252744 449074 252796 449080
rect 253216 447250 253244 452338
rect 253308 447914 253336 458866
rect 253296 447908 253348 447914
rect 253296 447850 253348 447856
rect 252664 447222 253152 447250
rect 253216 447222 253336 447250
rect 252744 446752 252796 446758
rect 252744 446694 252796 446700
rect 252756 443972 252784 446694
rect 252928 446276 252980 446282
rect 252928 446218 252980 446224
rect 252940 443972 252968 446218
rect 253124 443972 253152 447222
rect 253308 443972 253336 447222
rect 253480 444508 253532 444514
rect 253480 444450 253532 444456
rect 253492 443972 253520 444450
rect 253676 443972 253704 460906
rect 253848 449608 253900 449614
rect 253848 449550 253900 449556
rect 253860 443972 253888 449550
rect 253940 446412 253992 446418
rect 253940 446354 253992 446360
rect 253952 444802 253980 446354
rect 254044 445210 254072 460906
rect 254124 452600 254176 452606
rect 254124 452542 254176 452548
rect 254136 445398 254164 452542
rect 254584 452464 254636 452470
rect 254584 452406 254636 452412
rect 254124 445392 254176 445398
rect 254124 445334 254176 445340
rect 254044 445182 254256 445210
rect 253952 444774 254072 444802
rect 254044 443972 254072 444774
rect 254228 443972 254256 445182
rect 254400 444440 254452 444446
rect 254400 444382 254452 444388
rect 254412 443972 254440 444382
rect 254596 443972 254624 452406
rect 254768 450764 254820 450770
rect 254768 450706 254820 450712
rect 254780 443972 254808 450706
rect 254964 443972 254992 460906
rect 255872 452532 255924 452538
rect 255872 452474 255924 452480
rect 255688 450696 255740 450702
rect 255688 450638 255740 450644
rect 255320 450628 255372 450634
rect 255320 450570 255372 450576
rect 255332 448254 255360 450570
rect 255412 450560 255464 450566
rect 255412 450502 255464 450508
rect 255424 449585 255452 450502
rect 255410 449576 255466 449585
rect 255410 449511 255466 449520
rect 255412 448996 255464 449002
rect 255412 448938 255464 448944
rect 255320 448248 255372 448254
rect 255320 448190 255372 448196
rect 255424 446554 255452 448938
rect 255412 446548 255464 446554
rect 255412 446490 255464 446496
rect 255502 446448 255558 446457
rect 255502 446383 255558 446392
rect 255320 446344 255372 446350
rect 255320 446286 255372 446292
rect 255136 445392 255188 445398
rect 255136 445334 255188 445340
rect 255148 443972 255176 445334
rect 255332 443972 255360 446286
rect 255516 443972 255544 446383
rect 255700 443972 255728 450638
rect 255884 443972 255912 452474
rect 281000 452062 281028 596158
rect 281080 580508 281132 580514
rect 281080 580450 281132 580456
rect 280988 452056 281040 452062
rect 280988 451998 281040 452004
rect 256056 450832 256108 450838
rect 256056 450774 256108 450780
rect 256068 443972 256096 450774
rect 281092 449614 281120 580450
rect 281552 487966 281580 700266
rect 281632 596420 281684 596426
rect 281632 596362 281684 596368
rect 281540 487960 281592 487966
rect 281540 487902 281592 487908
rect 281644 452198 281672 596362
rect 282184 592680 282236 592686
rect 282184 592622 282236 592628
rect 281724 581664 281776 581670
rect 281724 581606 281776 581612
rect 281632 452192 281684 452198
rect 281632 452134 281684 452140
rect 281080 449608 281132 449614
rect 256422 449576 256478 449585
rect 281080 449550 281132 449556
rect 256422 449511 256478 449520
rect 256240 448248 256292 448254
rect 256240 448190 256292 448196
rect 256252 443972 256280 448190
rect 256332 446140 256384 446146
rect 256332 446082 256384 446088
rect 256344 443834 256372 446082
rect 256436 444145 256464 449511
rect 281736 449342 281764 581606
rect 282092 580576 282144 580582
rect 282092 580518 282144 580524
rect 281816 580440 281868 580446
rect 281816 580382 281868 580388
rect 281828 449546 281856 580382
rect 281908 580372 281960 580378
rect 281908 580314 281960 580320
rect 281816 449540 281868 449546
rect 281816 449482 281868 449488
rect 281920 449478 281948 580314
rect 282000 580304 282052 580310
rect 282000 580246 282052 580252
rect 281908 449472 281960 449478
rect 281908 449414 281960 449420
rect 282012 449410 282040 580246
rect 282104 452606 282132 580518
rect 282092 452600 282144 452606
rect 282092 452542 282144 452548
rect 282000 449404 282052 449410
rect 282000 449346 282052 449352
rect 281724 449336 281776 449342
rect 281724 449278 281776 449284
rect 258552 446962 258948 446978
rect 282196 446962 282224 592622
rect 282276 588600 282328 588606
rect 282276 588542 282328 588548
rect 282288 447098 282316 588542
rect 282368 580304 282420 580310
rect 282368 580246 282420 580252
rect 282276 447092 282328 447098
rect 282276 447034 282328 447040
rect 258540 446956 258960 446962
rect 258592 446950 258908 446956
rect 258540 446898 258592 446904
rect 258908 446898 258960 446904
rect 282184 446956 282236 446962
rect 282184 446898 282236 446904
rect 258816 446888 258868 446894
rect 258816 446830 258868 446836
rect 256606 446584 256662 446593
rect 256606 446519 256608 446528
rect 256660 446519 256662 446528
rect 256608 446490 256660 446496
rect 256516 446480 256568 446486
rect 256516 446422 256568 446428
rect 256528 446026 256556 446422
rect 258828 446214 258856 446830
rect 264978 446720 265034 446729
rect 264978 446655 265034 446664
rect 258816 446208 258868 446214
rect 258816 446150 258868 446156
rect 256528 445998 256648 446026
rect 256516 445868 256568 445874
rect 256516 445810 256568 445816
rect 256422 444136 256478 444145
rect 256422 444071 256478 444080
rect 256436 443972 256464 444071
rect 256528 443902 256556 445810
rect 256620 443972 256648 445998
rect 256790 445768 256846 445777
rect 256790 445703 256846 445712
rect 256804 443972 256832 445703
rect 256516 443896 256568 443902
rect 256516 443838 256568 443844
rect 254492 443828 254544 443834
rect 254492 443770 254544 443776
rect 256148 443828 256200 443834
rect 256148 443770 256200 443776
rect 256332 443828 256384 443834
rect 256332 443770 256384 443776
rect 249892 443760 249944 443766
rect 249892 443702 249944 443708
rect 229836 443692 229888 443698
rect 229836 443634 229888 443640
rect 234436 443692 234488 443698
rect 234436 443634 234488 443640
rect 239956 443692 240008 443698
rect 239956 443634 240008 443640
rect 242716 443692 242768 443698
rect 242716 443634 242768 443640
rect 248972 443692 249024 443698
rect 248972 443634 249024 443640
rect 220082 443391 220138 443400
rect 225236 443420 225288 443426
rect 217508 443362 217560 443368
rect 225788 443420 225840 443426
rect 225288 443380 225368 443408
rect 225236 443362 225288 443368
rect 225340 443292 225368 443380
rect 226340 443420 226392 443426
rect 225840 443380 225920 443408
rect 225788 443362 225840 443368
rect 225892 443292 225920 443380
rect 228180 443420 228232 443426
rect 226392 443380 226472 443408
rect 226340 443362 226392 443368
rect 226444 443292 226472 443380
rect 229468 443420 229520 443426
rect 228232 443380 228312 443408
rect 228180 443362 228232 443368
rect 228284 443292 228312 443380
rect 229848 443408 229876 443634
rect 234448 443494 234476 443634
rect 239036 443556 239088 443562
rect 239036 443498 239088 443504
rect 234436 443488 234488 443494
rect 234436 443430 234488 443436
rect 233700 443420 233752 443426
rect 229848 443380 229968 443408
rect 229468 443362 229520 443368
rect 229940 443292 229968 443380
rect 233620 443380 233700 443408
rect 233620 443292 233648 443380
rect 239048 443408 239076 443498
rect 239968 443426 239996 443634
rect 242728 443426 242756 443634
rect 242900 443556 242952 443562
rect 242820 443516 242900 443544
rect 242820 443428 242848 443516
rect 242900 443498 242952 443504
rect 254504 443426 254532 443770
rect 256160 443426 256188 443770
rect 233700 443362 233752 443368
rect 238956 443380 239076 443408
rect 239220 443420 239272 443426
rect 238956 443292 238984 443380
rect 239956 443420 240008 443426
rect 239272 443380 239352 443408
rect 239220 443362 239272 443368
rect 239324 443292 239352 443380
rect 239956 443362 240008 443368
rect 242716 443420 242768 443426
rect 242716 443362 242768 443368
rect 254492 443420 254544 443426
rect 254492 443362 254544 443368
rect 256148 443420 256200 443426
rect 256148 443362 256200 443368
rect 207754 398848 207810 398857
rect 207754 398783 207810 398792
rect 208032 398812 208084 398818
rect 207664 398744 207716 398750
rect 207664 398686 207716 398692
rect 207020 398608 207072 398614
rect 207020 398550 207072 398556
rect 203524 398472 203576 398478
rect 202142 398440 202198 398449
rect 203524 398414 203576 398420
rect 202142 398375 202198 398384
rect 201500 397316 201552 397322
rect 201500 397258 201552 397264
rect 200120 354612 200172 354618
rect 200120 354554 200172 354560
rect 199660 320136 199712 320142
rect 199660 320078 199712 320084
rect 199568 215280 199620 215286
rect 199568 215222 199620 215228
rect 199476 111784 199528 111790
rect 199476 111726 199528 111732
rect 199384 20664 199436 20670
rect 199384 20606 199436 20612
rect 200132 16574 200160 354554
rect 194612 16546 195192 16574
rect 200132 16546 200344 16574
rect 194414 6624 194470 6633
rect 194414 6559 194470 6568
rect 194428 480 194456 6559
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 198740 16176 198792 16182
rect 198740 16118 198792 16124
rect 197912 6520 197964 6526
rect 197912 6462 197964 6468
rect 196808 3732 196860 3738
rect 196808 3674 196860 3680
rect 196820 480 196848 3674
rect 197924 480 197952 6462
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 16118
rect 200316 480 200344 16546
rect 201512 3534 201540 397258
rect 202156 180130 202184 398375
rect 202880 392760 202932 392766
rect 202880 392702 202932 392708
rect 202144 180124 202196 180130
rect 202144 180066 202196 180072
rect 202892 16574 202920 392702
rect 202892 16546 203472 16574
rect 201592 5432 201644 5438
rect 201592 5374 201644 5380
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 201604 2802 201632 5374
rect 202696 3528 202748 3534
rect 202696 3470 202748 3476
rect 201512 2774 201632 2802
rect 201512 480 201540 2774
rect 202708 480 202736 3470
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203536 4826 203564 398414
rect 204904 398336 204956 398342
rect 204904 398278 204956 398284
rect 204916 398138 204944 398278
rect 204904 398132 204956 398138
rect 204904 398074 204956 398080
rect 206284 397860 206336 397866
rect 206284 397802 206336 397808
rect 203614 397760 203670 397769
rect 203614 397695 203670 397704
rect 203628 169046 203656 397695
rect 203616 169040 203668 169046
rect 203616 168982 203668 168988
rect 206296 86290 206324 397802
rect 206284 86284 206336 86290
rect 206284 86226 206336 86232
rect 206190 7984 206246 7993
rect 206190 7919 206246 7928
rect 203524 4820 203576 4826
rect 203524 4762 203576 4768
rect 205088 4820 205140 4826
rect 205088 4762 205140 4768
rect 205100 480 205128 4762
rect 206204 480 206232 7919
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 398550
rect 207676 4010 207704 398686
rect 207664 4004 207716 4010
rect 207664 3946 207716 3952
rect 207768 3466 207796 398783
rect 208032 398754 208084 398760
rect 210056 398812 210108 398818
rect 210056 398754 210108 398760
rect 210240 398812 210292 398818
rect 210240 398754 210292 398760
rect 207940 398676 207992 398682
rect 207940 398618 207992 398624
rect 207848 398540 207900 398546
rect 207848 398482 207900 398488
rect 207860 82142 207888 398482
rect 207952 178702 207980 398618
rect 208044 355434 208072 398754
rect 209228 398404 209280 398410
rect 209228 398346 209280 398352
rect 209044 397588 209096 397594
rect 209044 397530 209096 397536
rect 208398 392864 208454 392873
rect 208398 392799 208454 392808
rect 208032 355428 208084 355434
rect 208032 355370 208084 355376
rect 207940 178696 207992 178702
rect 207940 178638 207992 178644
rect 207848 82136 207900 82142
rect 207848 82078 207900 82084
rect 208412 16574 208440 392799
rect 208412 16546 208624 16574
rect 207756 3460 207808 3466
rect 207756 3402 207808 3408
rect 208596 480 208624 16546
rect 209056 6186 209084 397530
rect 209136 394392 209188 394398
rect 209136 394334 209188 394340
rect 209044 6180 209096 6186
rect 209044 6122 209096 6128
rect 209148 4078 209176 394334
rect 209240 338774 209268 398346
rect 209780 398132 209832 398138
rect 209780 398074 209832 398080
rect 209792 394466 209820 398074
rect 210068 398002 210096 398754
rect 210148 398676 210200 398682
rect 210148 398618 210200 398624
rect 210160 398070 210188 398618
rect 210252 398546 210280 398754
rect 210240 398540 210292 398546
rect 210240 398482 210292 398488
rect 210148 398064 210200 398070
rect 210148 398006 210200 398012
rect 210056 397996 210108 398002
rect 210056 397938 210108 397944
rect 210240 397792 210292 397798
rect 210240 397734 210292 397740
rect 210252 397526 210280 397734
rect 210240 397520 210292 397526
rect 210344 397497 210372 400044
rect 210240 397462 210292 397468
rect 210330 397488 210386 397497
rect 210330 397423 210386 397432
rect 210330 397080 210386 397089
rect 210330 397015 210386 397024
rect 210344 396817 210372 397015
rect 210330 396808 210386 396817
rect 210330 396743 210386 396752
rect 209872 396704 209924 396710
rect 210436 396658 210464 400044
rect 210528 396710 210556 400044
rect 209872 396646 209924 396652
rect 209780 394460 209832 394466
rect 209780 394402 209832 394408
rect 209780 393916 209832 393922
rect 209780 393858 209832 393864
rect 209228 338768 209280 338774
rect 209228 338710 209280 338716
rect 209136 4072 209188 4078
rect 209136 4014 209188 4020
rect 209792 480 209820 393858
rect 209884 9042 209912 396646
rect 209964 396636 210016 396642
rect 209964 396578 210016 396584
rect 210068 396630 210464 396658
rect 210516 396704 210568 396710
rect 210516 396646 210568 396652
rect 209976 9110 210004 396578
rect 209964 9104 210016 9110
rect 209964 9046 210016 9052
rect 209872 9036 209924 9042
rect 209872 8978 209924 8984
rect 210068 8974 210096 396630
rect 210620 396522 210648 400044
rect 210712 398138 210740 400044
rect 210700 398132 210752 398138
rect 210700 398074 210752 398080
rect 210698 398032 210754 398041
rect 210698 397967 210754 397976
rect 210712 397769 210740 397967
rect 210698 397760 210754 397769
rect 210698 397695 210754 397704
rect 210804 397594 210832 400044
rect 210792 397588 210844 397594
rect 210792 397530 210844 397536
rect 210700 397520 210752 397526
rect 210700 397462 210752 397468
rect 210160 396494 210648 396522
rect 210160 13122 210188 396494
rect 210240 396432 210292 396438
rect 210240 396374 210292 396380
rect 210252 13190 210280 396374
rect 210332 396364 210384 396370
rect 210332 396306 210384 396312
rect 210344 177342 210372 396306
rect 210516 396160 210568 396166
rect 210516 396102 210568 396108
rect 210424 393984 210476 393990
rect 210424 393926 210476 393932
rect 210332 177336 210384 177342
rect 210332 177278 210384 177284
rect 210240 13184 210292 13190
rect 210240 13126 210292 13132
rect 210148 13116 210200 13122
rect 210148 13058 210200 13064
rect 210056 8968 210108 8974
rect 210056 8910 210108 8916
rect 210436 3738 210464 393926
rect 210528 393922 210556 396102
rect 210516 393916 210568 393922
rect 210516 393858 210568 393864
rect 210712 393802 210740 397462
rect 210792 397452 210844 397458
rect 210792 397394 210844 397400
rect 210528 393774 210740 393802
rect 210528 15978 210556 393774
rect 210804 393314 210832 397394
rect 210896 396642 210924 400044
rect 210884 396636 210936 396642
rect 210884 396578 210936 396584
rect 210988 396438 211016 400044
rect 210976 396432 211028 396438
rect 210976 396374 211028 396380
rect 211080 396370 211108 400044
rect 211172 398313 211200 400044
rect 211158 398304 211214 398313
rect 211158 398239 211214 398248
rect 211160 397520 211212 397526
rect 211160 397462 211212 397468
rect 211068 396364 211120 396370
rect 211068 396306 211120 396312
rect 210620 393286 210832 393314
rect 210620 352578 210648 393286
rect 210608 352572 210660 352578
rect 210608 352514 210660 352520
rect 210516 15972 210568 15978
rect 210516 15914 210568 15920
rect 211172 14754 211200 397462
rect 211264 396817 211292 400044
rect 211356 397497 211384 400044
rect 211448 397633 211476 400044
rect 211540 398585 211568 400044
rect 211526 398576 211582 398585
rect 211526 398511 211582 398520
rect 211528 397928 211580 397934
rect 211528 397870 211580 397876
rect 211434 397624 211490 397633
rect 211540 397594 211568 397870
rect 211632 397769 211660 400044
rect 211618 397760 211674 397769
rect 211618 397695 211674 397704
rect 211434 397559 211490 397568
rect 211528 397588 211580 397594
rect 211528 397530 211580 397536
rect 211342 397488 211398 397497
rect 211342 397423 211398 397432
rect 211620 397384 211672 397390
rect 211620 397326 211672 397332
rect 211632 396846 211660 397326
rect 211620 396840 211672 396846
rect 211250 396808 211306 396817
rect 211620 396782 211672 396788
rect 211250 396743 211306 396752
rect 211344 396704 211396 396710
rect 211724 396658 211752 400044
rect 211816 398478 211844 400044
rect 211804 398472 211856 398478
rect 211804 398414 211856 398420
rect 211908 397905 211936 400044
rect 211894 397896 211950 397905
rect 211894 397831 211950 397840
rect 211802 397624 211858 397633
rect 211802 397559 211858 397568
rect 211896 397588 211948 397594
rect 211344 396646 211396 396652
rect 211252 396636 211304 396642
rect 211252 396578 211304 396584
rect 211160 14748 211212 14754
rect 211160 14690 211212 14696
rect 211264 11762 211292 396578
rect 211356 14550 211384 396646
rect 211448 396630 211752 396658
rect 211344 14544 211396 14550
rect 211344 14486 211396 14492
rect 211448 14482 211476 396630
rect 211528 396568 211580 396574
rect 211528 396510 211580 396516
rect 211436 14476 211488 14482
rect 211436 14418 211488 14424
rect 211540 11830 211568 396510
rect 211816 14618 211844 397559
rect 211896 397530 211948 397536
rect 211908 15910 211936 397530
rect 212000 396642 212028 400044
rect 212092 396710 212120 400044
rect 212184 398410 212212 400044
rect 212172 398404 212224 398410
rect 212172 398346 212224 398352
rect 212276 398342 212304 400044
rect 212264 398336 212316 398342
rect 212170 398304 212226 398313
rect 212264 398278 212316 398284
rect 212170 398239 212226 398248
rect 212080 396704 212132 396710
rect 212080 396646 212132 396652
rect 211988 396636 212040 396642
rect 211988 396578 212040 396584
rect 212184 395350 212212 398239
rect 212262 397896 212318 397905
rect 212262 397831 212318 397840
rect 212172 395344 212224 395350
rect 212172 395286 212224 395292
rect 212276 393314 212304 397831
rect 212368 396574 212396 400044
rect 212460 398313 212488 400044
rect 212446 398304 212502 398313
rect 212446 398239 212502 398248
rect 212448 398132 212500 398138
rect 212448 398074 212500 398080
rect 212356 396568 212408 396574
rect 212356 396510 212408 396516
rect 212460 394330 212488 398074
rect 212552 397769 212580 400044
rect 212538 397760 212594 397769
rect 212538 397695 212594 397704
rect 212644 397497 212672 400044
rect 212630 397488 212686 397497
rect 212630 397423 212686 397432
rect 212540 397248 212592 397254
rect 212540 397190 212592 397196
rect 212552 396778 212580 397190
rect 212736 396930 212764 400044
rect 212828 398041 212856 400044
rect 212814 398032 212870 398041
rect 212814 397967 212870 397976
rect 212644 396902 212764 396930
rect 212540 396772 212592 396778
rect 212540 396714 212592 396720
rect 212644 396658 212672 396902
rect 212724 396840 212776 396846
rect 212724 396782 212776 396788
rect 212552 396630 212672 396658
rect 212552 395418 212580 396630
rect 212632 396500 212684 396506
rect 212632 396442 212684 396448
rect 212540 395412 212592 395418
rect 212540 395354 212592 395360
rect 212448 394324 212500 394330
rect 212448 394266 212500 394272
rect 212092 393286 212304 393314
rect 212092 354210 212120 393286
rect 212080 354204 212132 354210
rect 212080 354146 212132 354152
rect 211896 15904 211948 15910
rect 211896 15846 211948 15852
rect 211804 14612 211856 14618
rect 211804 14554 211856 14560
rect 212644 12034 212672 396442
rect 212632 12028 212684 12034
rect 212632 11970 212684 11976
rect 212736 11966 212764 396782
rect 212920 396778 212948 400044
rect 213012 397633 213040 400044
rect 212998 397624 213054 397633
rect 212998 397559 213054 397568
rect 212908 396772 212960 396778
rect 212908 396714 212960 396720
rect 212816 396704 212868 396710
rect 212816 396646 212868 396652
rect 212828 14822 212856 396646
rect 212908 396636 212960 396642
rect 212908 396578 212960 396584
rect 212816 14816 212868 14822
rect 212816 14758 212868 14764
rect 212920 14686 212948 396578
rect 213000 396568 213052 396574
rect 213000 396510 213052 396516
rect 213012 354074 213040 396510
rect 213000 354068 213052 354074
rect 213000 354010 213052 354016
rect 213104 354006 213132 400044
rect 213196 396846 213224 400044
rect 213184 396840 213236 396846
rect 213184 396782 213236 396788
rect 213288 396642 213316 400044
rect 213380 398449 213408 400044
rect 213366 398440 213422 398449
rect 213366 398375 213422 398384
rect 213368 398336 213420 398342
rect 213368 398278 213420 398284
rect 213380 396930 213408 398278
rect 213472 397254 213500 400044
rect 213564 397526 213592 400044
rect 213552 397520 213604 397526
rect 213552 397462 213604 397468
rect 213460 397248 213512 397254
rect 213460 397190 213512 397196
rect 213380 396902 213500 396930
rect 213368 396772 213420 396778
rect 213368 396714 213420 396720
rect 213276 396636 213328 396642
rect 213276 396578 213328 396584
rect 213184 395956 213236 395962
rect 213184 395898 213236 395904
rect 213092 354000 213144 354006
rect 213092 353942 213144 353948
rect 212908 14680 212960 14686
rect 212908 14622 212960 14628
rect 212724 11960 212776 11966
rect 212724 11902 212776 11908
rect 211528 11824 211580 11830
rect 211528 11766 211580 11772
rect 211252 11756 211304 11762
rect 211252 11698 211304 11704
rect 210976 4072 211028 4078
rect 210976 4014 211028 4020
rect 210424 3732 210476 3738
rect 210424 3674 210476 3680
rect 210988 480 211016 4014
rect 213196 3942 213224 395898
rect 213274 394768 213330 394777
rect 213274 394703 213330 394712
rect 213184 3936 213236 3942
rect 213184 3878 213236 3884
rect 213288 3806 213316 394703
rect 213380 11898 213408 396714
rect 213472 395962 213500 396902
rect 213656 396574 213684 400044
rect 213644 396568 213696 396574
rect 213644 396510 213696 396516
rect 213748 396506 213776 400044
rect 213840 396710 213868 400044
rect 213828 396704 213880 396710
rect 213828 396646 213880 396652
rect 213736 396500 213788 396506
rect 213736 396442 213788 396448
rect 213460 395956 213512 395962
rect 213460 395898 213512 395904
rect 213932 395457 213960 400044
rect 214024 398857 214052 400044
rect 214010 398848 214066 398857
rect 214010 398783 214066 398792
rect 214012 398676 214064 398682
rect 214012 398618 214064 398624
rect 214024 395962 214052 398618
rect 214116 397497 214144 400044
rect 214208 397769 214236 400044
rect 214194 397760 214250 397769
rect 214194 397695 214250 397704
rect 214300 397633 214328 400044
rect 214286 397624 214342 397633
rect 214286 397559 214342 397568
rect 214102 397488 214158 397497
rect 214102 397423 214158 397432
rect 214392 396930 214420 400044
rect 214484 398682 214512 400044
rect 214472 398676 214524 398682
rect 214472 398618 214524 398624
rect 214300 396902 214420 396930
rect 214104 396772 214156 396778
rect 214104 396714 214156 396720
rect 214012 395956 214064 395962
rect 214012 395898 214064 395904
rect 214012 395820 214064 395826
rect 214012 395762 214064 395768
rect 213918 395448 213974 395457
rect 213918 395383 213974 395392
rect 213368 11892 213420 11898
rect 213368 11834 213420 11840
rect 214024 9246 214052 395762
rect 214012 9240 214064 9246
rect 214012 9182 214064 9188
rect 214116 9178 214144 396714
rect 214196 396704 214248 396710
rect 214196 396646 214248 396652
rect 214208 13394 214236 396646
rect 214196 13388 214248 13394
rect 214196 13330 214248 13336
rect 214300 13258 214328 396902
rect 214576 396778 214604 400044
rect 214564 396772 214616 396778
rect 214564 396714 214616 396720
rect 214472 396636 214524 396642
rect 214472 396578 214524 396584
rect 214380 395956 214432 395962
rect 214380 395898 214432 395904
rect 214392 395486 214420 395898
rect 214380 395480 214432 395486
rect 214380 395422 214432 395428
rect 214380 395208 214432 395214
rect 214380 395150 214432 395156
rect 214392 13326 214420 395150
rect 214484 14890 214512 396578
rect 214564 396568 214616 396574
rect 214564 396510 214616 396516
rect 214576 354142 214604 396510
rect 214668 395214 214696 400044
rect 214760 396642 214788 400044
rect 214748 396636 214800 396642
rect 214748 396578 214800 396584
rect 214852 395826 214880 400044
rect 214944 396710 214972 400044
rect 215036 397594 215064 400044
rect 215024 397588 215076 397594
rect 215024 397530 215076 397536
rect 215024 397452 215076 397458
rect 215024 397394 215076 397400
rect 214932 396704 214984 396710
rect 214932 396646 214984 396652
rect 214840 395820 214892 395826
rect 214840 395762 214892 395768
rect 214656 395208 214708 395214
rect 214656 395150 214708 395156
rect 215036 395026 215064 397394
rect 214668 394998 215064 395026
rect 214668 392630 214696 394998
rect 215128 393314 215156 400044
rect 215220 396574 215248 400044
rect 215312 397497 215340 400044
rect 215298 397488 215354 397497
rect 215298 397423 215354 397432
rect 215404 397089 215432 400044
rect 215496 397633 215524 400044
rect 215588 397769 215616 400044
rect 215574 397760 215630 397769
rect 215574 397695 215630 397704
rect 215482 397624 215538 397633
rect 215482 397559 215538 397568
rect 215390 397080 215446 397089
rect 215390 397015 215446 397024
rect 215208 396568 215260 396574
rect 215208 396510 215260 396516
rect 215300 394664 215352 394670
rect 215300 394606 215352 394612
rect 215312 394194 215340 394606
rect 215392 394596 215444 394602
rect 215392 394538 215444 394544
rect 215300 394188 215352 394194
rect 215300 394130 215352 394136
rect 214760 393286 215156 393314
rect 214656 392624 214708 392630
rect 214656 392566 214708 392572
rect 214564 354136 214616 354142
rect 214564 354078 214616 354084
rect 214472 14884 214524 14890
rect 214472 14826 214524 14832
rect 214380 13320 214432 13326
rect 214380 13262 214432 13268
rect 214288 13252 214340 13258
rect 214288 13194 214340 13200
rect 214760 9314 214788 393286
rect 215404 9450 215432 394538
rect 215576 394188 215628 394194
rect 215576 394130 215628 394136
rect 215484 393780 215536 393786
rect 215484 393722 215536 393728
rect 215496 10470 215524 393722
rect 215484 10464 215536 10470
rect 215484 10406 215536 10412
rect 215588 10402 215616 394130
rect 215680 394058 215708 400044
rect 215668 394052 215720 394058
rect 215668 393994 215720 394000
rect 215668 393916 215720 393922
rect 215668 393858 215720 393864
rect 215680 13598 215708 393858
rect 215772 393666 215800 400044
rect 215864 397905 215892 400044
rect 215850 397896 215906 397905
rect 215850 397831 215906 397840
rect 215956 394602 215984 400044
rect 215944 394596 215996 394602
rect 215944 394538 215996 394544
rect 216048 393938 216076 400044
rect 215956 393910 216076 393938
rect 215956 393825 215984 393910
rect 216036 393848 216088 393854
rect 215942 393816 215998 393825
rect 216036 393790 216088 393796
rect 215942 393751 215998 393760
rect 215944 393712 215996 393718
rect 215772 393638 215892 393666
rect 215944 393654 215996 393660
rect 215758 393544 215814 393553
rect 215758 393479 215814 393488
rect 215668 13592 215720 13598
rect 215668 13534 215720 13540
rect 215772 13530 215800 393479
rect 215760 13524 215812 13530
rect 215760 13466 215812 13472
rect 215864 13462 215892 393638
rect 215852 13456 215904 13462
rect 215852 13398 215904 13404
rect 215576 10396 215628 10402
rect 215576 10338 215628 10344
rect 215392 9444 215444 9450
rect 215392 9386 215444 9392
rect 214748 9308 214800 9314
rect 214748 9250 214800 9256
rect 214104 9172 214156 9178
rect 214104 9114 214156 9120
rect 213368 4004 213420 4010
rect 213368 3946 213420 3952
rect 213276 3800 213328 3806
rect 213276 3742 213328 3748
rect 212172 3732 212224 3738
rect 212172 3674 212224 3680
rect 212184 480 212212 3674
rect 213380 480 213408 3946
rect 215668 3936 215720 3942
rect 215668 3878 215720 3884
rect 214472 3800 214524 3806
rect 214472 3742 214524 3748
rect 214484 480 214512 3742
rect 215680 480 215708 3878
rect 215956 3874 215984 393654
rect 216048 177410 216076 393790
rect 216140 351218 216168 400044
rect 216232 394194 216260 400044
rect 216220 394188 216272 394194
rect 216220 394130 216272 394136
rect 216220 394052 216272 394058
rect 216220 393994 216272 394000
rect 216128 351212 216180 351218
rect 216128 351154 216180 351160
rect 216036 177404 216088 177410
rect 216036 177346 216088 177352
rect 216232 9382 216260 393994
rect 216324 393922 216352 400044
rect 216416 395554 216444 400044
rect 216404 395548 216456 395554
rect 216404 395490 216456 395496
rect 216404 394732 216456 394738
rect 216404 394674 216456 394680
rect 216312 393916 216364 393922
rect 216312 393858 216364 393864
rect 216416 393718 216444 394674
rect 216508 393786 216536 400044
rect 216600 393854 216628 400044
rect 216692 397633 216720 400044
rect 216678 397624 216734 397633
rect 216678 397559 216734 397568
rect 216784 397497 216812 400044
rect 216876 397769 216904 400044
rect 216968 399090 216996 400044
rect 216956 399084 217008 399090
rect 216956 399026 217008 399032
rect 216954 398712 217010 398721
rect 216954 398647 217010 398656
rect 216968 397798 216996 398647
rect 217060 397905 217088 400044
rect 217046 397896 217102 397905
rect 217046 397831 217102 397840
rect 216956 397792 217008 397798
rect 216862 397760 216918 397769
rect 216956 397734 217008 397740
rect 217048 397792 217100 397798
rect 217048 397734 217100 397740
rect 216862 397695 216918 397704
rect 216770 397488 216826 397497
rect 216770 397423 216826 397432
rect 216956 394188 217008 394194
rect 216956 394130 217008 394136
rect 216864 394052 216916 394058
rect 216864 393994 216916 394000
rect 216588 393848 216640 393854
rect 216588 393790 216640 393796
rect 216496 393780 216548 393786
rect 216496 393722 216548 393728
rect 216404 393712 216456 393718
rect 216404 393654 216456 393660
rect 216876 10674 216904 393994
rect 216968 354346 216996 394130
rect 217060 392698 217088 397734
rect 217048 392692 217100 392698
rect 217048 392634 217100 392640
rect 217152 392306 217180 400044
rect 217244 399226 217272 400044
rect 217232 399220 217284 399226
rect 217232 399162 217284 399168
rect 217232 399084 217284 399090
rect 217232 399026 217284 399032
rect 217244 398857 217272 399026
rect 217230 398848 217286 398857
rect 217230 398783 217286 398792
rect 217232 398676 217284 398682
rect 217232 398618 217284 398624
rect 217244 397934 217272 398618
rect 217232 397928 217284 397934
rect 217232 397870 217284 397876
rect 217232 397452 217284 397458
rect 217232 397394 217284 397400
rect 217244 396166 217272 397394
rect 217232 396160 217284 396166
rect 217232 396102 217284 396108
rect 217060 392278 217180 392306
rect 216956 354340 217008 354346
rect 216956 354282 217008 354288
rect 217060 354278 217088 392278
rect 217140 392216 217192 392222
rect 217140 392158 217192 392164
rect 217152 354414 217180 392158
rect 217336 389298 217364 400044
rect 217428 394194 217456 400044
rect 217520 398857 217548 400044
rect 217612 399022 217640 400044
rect 217600 399016 217652 399022
rect 217600 398958 217652 398964
rect 217704 398954 217732 400044
rect 217692 398948 217744 398954
rect 217692 398890 217744 398896
rect 217506 398848 217562 398857
rect 217506 398783 217562 398792
rect 217690 398848 217746 398857
rect 217690 398783 217746 398792
rect 217508 398744 217560 398750
rect 217508 398686 217560 398692
rect 217600 398744 217652 398750
rect 217600 398686 217652 398692
rect 217520 395690 217548 398686
rect 217508 395684 217560 395690
rect 217508 395626 217560 395632
rect 217416 394188 217468 394194
rect 217416 394130 217468 394136
rect 217612 389314 217640 398686
rect 217704 394126 217732 398783
rect 217796 398682 217824 400044
rect 217784 398676 217836 398682
rect 217784 398618 217836 398624
rect 217784 398540 217836 398546
rect 217784 398482 217836 398488
rect 217796 397798 217824 398482
rect 217784 397792 217836 397798
rect 217784 397734 217836 397740
rect 217784 397656 217836 397662
rect 217784 397598 217836 397604
rect 217796 396982 217824 397598
rect 217784 396976 217836 396982
rect 217784 396918 217836 396924
rect 217692 394120 217744 394126
rect 217692 394062 217744 394068
rect 217888 394058 217916 400044
rect 217876 394052 217928 394058
rect 217876 393994 217928 394000
rect 217980 392222 218008 400044
rect 218072 397633 218100 400044
rect 218058 397624 218114 397633
rect 218058 397559 218114 397568
rect 218164 397497 218192 400044
rect 218256 397769 218284 400044
rect 218348 398070 218376 400044
rect 218336 398064 218388 398070
rect 218336 398006 218388 398012
rect 218242 397760 218298 397769
rect 218242 397695 218298 397704
rect 218150 397488 218206 397497
rect 218150 397423 218206 397432
rect 218244 394120 218296 394126
rect 218244 394062 218296 394068
rect 217968 392216 218020 392222
rect 217968 392158 218020 392164
rect 217324 389292 217376 389298
rect 217324 389234 217376 389240
rect 217428 389286 217640 389314
rect 217428 386414 217456 389286
rect 217508 389088 217560 389094
rect 217508 389030 217560 389036
rect 217244 386386 217456 386414
rect 217140 354408 217192 354414
rect 217140 354350 217192 354356
rect 217048 354272 217100 354278
rect 217048 354214 217100 354220
rect 216956 89004 217008 89010
rect 216956 88946 217008 88952
rect 216864 10668 216916 10674
rect 216864 10610 216916 10616
rect 216220 9376 216272 9382
rect 216220 9318 216272 9324
rect 216968 6914 216996 88946
rect 217244 10606 217272 386386
rect 217232 10600 217284 10606
rect 217232 10542 217284 10548
rect 217520 10538 217548 389030
rect 218256 12102 218284 394062
rect 218440 393922 218468 400044
rect 218428 393916 218480 393922
rect 218428 393858 218480 393864
rect 218336 393848 218388 393854
rect 218336 393790 218388 393796
rect 218348 12170 218376 393790
rect 218428 393780 218480 393786
rect 218428 393722 218480 393728
rect 218440 16046 218468 393722
rect 218532 355366 218560 400044
rect 218624 397390 218652 400044
rect 218612 397384 218664 397390
rect 218612 397326 218664 397332
rect 218612 394052 218664 394058
rect 218716 394040 218744 400044
rect 218808 397594 218836 400044
rect 218900 398002 218928 400044
rect 218888 397996 218940 398002
rect 218888 397938 218940 397944
rect 218796 397588 218848 397594
rect 218796 397530 218848 397536
rect 218888 397588 218940 397594
rect 218888 397530 218940 397536
rect 218900 394670 218928 397530
rect 218888 394664 218940 394670
rect 218888 394606 218940 394612
rect 218992 394126 219020 400044
rect 218980 394120 219032 394126
rect 218980 394062 219032 394068
rect 219084 394058 219112 400044
rect 219072 394052 219124 394058
rect 218716 394012 218928 394040
rect 218612 393994 218664 394000
rect 218520 355360 218572 355366
rect 218520 355302 218572 355308
rect 218520 351212 218572 351218
rect 218520 351154 218572 351160
rect 218428 16040 218480 16046
rect 218428 15982 218480 15988
rect 218336 12164 218388 12170
rect 218336 12106 218388 12112
rect 218244 12096 218296 12102
rect 218244 12038 218296 12044
rect 217508 10532 217560 10538
rect 217508 10474 217560 10480
rect 218532 6914 218560 351154
rect 218624 177478 218652 393994
rect 218796 393916 218848 393922
rect 218796 393858 218848 393864
rect 218612 177472 218664 177478
rect 218612 177414 218664 177420
rect 218808 10742 218836 393858
rect 218900 389174 218928 394012
rect 219072 393994 219124 394000
rect 219176 393786 219204 400044
rect 219268 393854 219296 400044
rect 219360 399129 219388 400044
rect 219346 399120 219402 399129
rect 219346 399055 219402 399064
rect 219452 399022 219480 400044
rect 219348 399016 219400 399022
rect 219348 398958 219400 398964
rect 219440 399016 219492 399022
rect 219440 398958 219492 398964
rect 219360 398834 219388 398958
rect 219360 398806 219480 398834
rect 219346 398712 219402 398721
rect 219346 398647 219402 398656
rect 219360 395622 219388 398647
rect 219452 397934 219480 398806
rect 219440 397928 219492 397934
rect 219440 397870 219492 397876
rect 219440 397792 219492 397798
rect 219440 397734 219492 397740
rect 219348 395616 219400 395622
rect 219348 395558 219400 395564
rect 219256 393848 219308 393854
rect 219256 393790 219308 393796
rect 219164 393780 219216 393786
rect 219164 393722 219216 393728
rect 218900 389146 219020 389174
rect 218992 10810 219020 389146
rect 218980 10804 219032 10810
rect 218980 10746 219032 10752
rect 218796 10736 218848 10742
rect 218796 10678 218848 10684
rect 216876 6886 216996 6914
rect 218072 6886 218560 6914
rect 215944 3868 215996 3874
rect 215944 3810 215996 3816
rect 216876 480 216904 6886
rect 218072 480 218100 6886
rect 219256 3868 219308 3874
rect 219256 3810 219308 3816
rect 219268 480 219296 3810
rect 219452 490 219480 397734
rect 219544 397497 219572 400044
rect 219530 397488 219586 397497
rect 219530 397423 219586 397432
rect 219636 395729 219664 400044
rect 219728 397497 219756 400044
rect 219820 397633 219848 400044
rect 219806 397624 219862 397633
rect 219806 397559 219862 397568
rect 219714 397488 219770 397497
rect 219714 397423 219770 397432
rect 219622 395720 219678 395729
rect 219622 395655 219678 395664
rect 219532 394120 219584 394126
rect 219532 394062 219584 394068
rect 219544 3602 219572 394062
rect 219808 394052 219860 394058
rect 219808 393994 219860 394000
rect 219716 393916 219768 393922
rect 219716 393858 219768 393864
rect 219624 393848 219676 393854
rect 219624 393790 219676 393796
rect 219636 3670 219664 393790
rect 219728 4894 219756 393858
rect 219820 6254 219848 393994
rect 219912 16114 219940 400044
rect 220004 177546 220032 400044
rect 220096 398206 220124 400044
rect 220084 398200 220136 398206
rect 220084 398142 220136 398148
rect 220084 397520 220136 397526
rect 220084 397462 220136 397468
rect 219992 177540 220044 177546
rect 219992 177482 220044 177488
rect 219900 16108 219952 16114
rect 219900 16050 219952 16056
rect 220096 7886 220124 397462
rect 220188 393922 220216 400044
rect 220280 394058 220308 400044
rect 220372 394126 220400 400044
rect 220464 394262 220492 400044
rect 220556 396914 220584 400044
rect 220544 396908 220596 396914
rect 220544 396850 220596 396856
rect 220452 394256 220504 394262
rect 220452 394198 220504 394204
rect 220360 394120 220412 394126
rect 220360 394062 220412 394068
rect 220268 394052 220320 394058
rect 220268 393994 220320 394000
rect 220176 393916 220228 393922
rect 220176 393858 220228 393864
rect 220648 393854 220676 400044
rect 220740 397594 220768 400044
rect 220832 397662 220860 400044
rect 220924 397769 220952 400044
rect 220910 397760 220966 397769
rect 220910 397695 220966 397704
rect 220820 397656 220872 397662
rect 221016 397633 221044 400044
rect 220820 397598 220872 397604
rect 221002 397624 221058 397633
rect 220728 397588 220780 397594
rect 221002 397559 221058 397568
rect 220728 397530 220780 397536
rect 221108 397497 221136 400044
rect 221200 397633 221228 400044
rect 221186 397624 221242 397633
rect 221186 397559 221242 397568
rect 221094 397488 221150 397497
rect 221094 397423 221150 397432
rect 221096 394324 221148 394330
rect 221096 394266 221148 394272
rect 220912 394188 220964 394194
rect 220912 394130 220964 394136
rect 220636 393848 220688 393854
rect 220636 393790 220688 393796
rect 220820 351960 220872 351966
rect 220820 351902 220872 351908
rect 220832 11762 220860 351902
rect 220820 11756 220872 11762
rect 220820 11698 220872 11704
rect 220084 7880 220136 7886
rect 220084 7822 220136 7828
rect 219808 6248 219860 6254
rect 219808 6190 219860 6196
rect 220924 5030 220952 394130
rect 221004 393848 221056 393854
rect 221004 393790 221056 393796
rect 221016 7818 221044 393790
rect 221004 7812 221056 7818
rect 221004 7754 221056 7760
rect 221108 7682 221136 394266
rect 221188 394120 221240 394126
rect 221188 394062 221240 394068
rect 221200 7750 221228 394062
rect 221188 7744 221240 7750
rect 221188 7686 221240 7692
rect 221096 7676 221148 7682
rect 221096 7618 221148 7624
rect 221292 7614 221320 400044
rect 221384 394040 221412 400044
rect 221476 394210 221504 400044
rect 221568 394330 221596 400044
rect 221660 397050 221688 400044
rect 221648 397044 221700 397050
rect 221648 396986 221700 396992
rect 221556 394324 221608 394330
rect 221556 394266 221608 394272
rect 221476 394182 221688 394210
rect 221556 394052 221608 394058
rect 221384 394012 221504 394040
rect 221372 393916 221424 393922
rect 221372 393858 221424 393864
rect 221384 46238 221412 393858
rect 221476 351286 221504 394012
rect 221556 393994 221608 394000
rect 221568 352646 221596 393994
rect 221556 352640 221608 352646
rect 221556 352582 221608 352588
rect 221464 351280 221516 351286
rect 221464 351222 221516 351228
rect 221372 46232 221424 46238
rect 221372 46174 221424 46180
rect 221372 11756 221424 11762
rect 221372 11698 221424 11704
rect 221280 7608 221332 7614
rect 221280 7550 221332 7556
rect 220912 5024 220964 5030
rect 220912 4966 220964 4972
rect 219716 4888 219768 4894
rect 219716 4830 219768 4836
rect 219624 3664 219676 3670
rect 219624 3606 219676 3612
rect 219532 3596 219584 3602
rect 219532 3538 219584 3544
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 219452 462 220032 490
rect 220004 354 220032 462
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221384 354 221412 11698
rect 221660 4962 221688 394182
rect 221752 393922 221780 400044
rect 221844 394126 221872 400044
rect 221832 394120 221884 394126
rect 221832 394062 221884 394068
rect 221936 394058 221964 400044
rect 222028 394194 222056 400044
rect 222016 394188 222068 394194
rect 222016 394130 222068 394136
rect 221924 394052 221976 394058
rect 221924 393994 221976 394000
rect 221740 393916 221792 393922
rect 221740 393858 221792 393864
rect 222120 393854 222148 400044
rect 222212 397769 222240 400044
rect 222198 397760 222254 397769
rect 222198 397695 222254 397704
rect 222200 397656 222252 397662
rect 222200 397598 222252 397604
rect 222108 393848 222160 393854
rect 222108 393790 222160 393796
rect 222212 16574 222240 397598
rect 222304 397497 222332 400044
rect 222396 397526 222424 400044
rect 222384 397520 222436 397526
rect 222290 397488 222346 397497
rect 222384 397462 222436 397468
rect 222290 397423 222346 397432
rect 222384 394188 222436 394194
rect 222384 394130 222436 394136
rect 222212 16546 222332 16574
rect 221648 4956 221700 4962
rect 221648 4898 221700 4904
rect 222304 3482 222332 16546
rect 222396 5166 222424 394130
rect 222488 393922 222516 400044
rect 222476 393916 222528 393922
rect 222476 393858 222528 393864
rect 222580 389450 222608 400044
rect 222488 389422 222608 389450
rect 222384 5160 222436 5166
rect 222384 5102 222436 5108
rect 222488 5098 222516 389422
rect 222568 389360 222620 389366
rect 222568 389302 222620 389308
rect 222580 5302 222608 389302
rect 222672 7954 222700 400044
rect 222764 397118 222792 400044
rect 222856 398546 222884 400044
rect 222844 398540 222896 398546
rect 222844 398482 222896 398488
rect 222752 397112 222804 397118
rect 222752 397054 222804 397060
rect 222752 396364 222804 396370
rect 222752 396306 222804 396312
rect 222764 392714 222792 396306
rect 222948 394194 222976 400044
rect 222936 394188 222988 394194
rect 222936 394130 222988 394136
rect 222936 393916 222988 393922
rect 222936 393858 222988 393864
rect 222764 392686 222884 392714
rect 222752 391060 222804 391066
rect 222752 391002 222804 391008
rect 222764 46306 222792 391002
rect 222752 46300 222804 46306
rect 222752 46242 222804 46248
rect 222660 7948 222712 7954
rect 222660 7890 222712 7896
rect 222568 5296 222620 5302
rect 222568 5238 222620 5244
rect 222476 5092 222528 5098
rect 222476 5034 222528 5040
rect 222856 3874 222884 392686
rect 222948 177614 222976 393858
rect 223040 391066 223068 400044
rect 223132 398342 223160 400044
rect 223120 398336 223172 398342
rect 223120 398278 223172 398284
rect 223028 391060 223080 391066
rect 223028 391002 223080 391008
rect 223224 389174 223252 400044
rect 223316 394738 223344 400044
rect 223408 398478 223436 400044
rect 223396 398472 223448 398478
rect 223396 398414 223448 398420
rect 223304 394732 223356 394738
rect 223304 394674 223356 394680
rect 223500 389366 223528 400044
rect 223592 397769 223620 400044
rect 223684 398274 223712 400044
rect 223672 398268 223724 398274
rect 223672 398210 223724 398216
rect 223578 397760 223634 397769
rect 223578 397695 223634 397704
rect 223776 397497 223804 400044
rect 223868 397633 223896 400044
rect 223854 397624 223910 397633
rect 223854 397559 223910 397568
rect 223960 397497 223988 400044
rect 223762 397488 223818 397497
rect 223762 397423 223818 397432
rect 223946 397488 224002 397497
rect 223946 397423 224002 397432
rect 223764 394324 223816 394330
rect 223764 394266 223816 394272
rect 223488 389360 223540 389366
rect 223488 389302 223540 389308
rect 223224 389146 223528 389174
rect 222936 177608 222988 177614
rect 222936 177550 222988 177556
rect 223500 5234 223528 389146
rect 223776 6322 223804 394266
rect 223856 394188 223908 394194
rect 223856 394130 223908 394136
rect 223868 6390 223896 394130
rect 223948 394120 224000 394126
rect 223948 394062 224000 394068
rect 223960 6458 223988 394062
rect 224052 393922 224080 400044
rect 224040 393916 224092 393922
rect 224040 393858 224092 393864
rect 224144 392306 224172 400044
rect 224236 394398 224264 400044
rect 224224 394392 224276 394398
rect 224224 394334 224276 394340
rect 224328 394330 224356 400044
rect 224316 394324 224368 394330
rect 224316 394266 224368 394272
rect 224420 394210 224448 400044
rect 224512 394534 224540 400044
rect 224500 394528 224552 394534
rect 224500 394470 224552 394476
rect 224052 392278 224172 392306
rect 224236 394182 224448 394210
rect 224604 394194 224632 400044
rect 224592 394188 224644 394194
rect 224052 354482 224080 392278
rect 224236 392170 224264 394182
rect 224592 394130 224644 394136
rect 224316 394052 224368 394058
rect 224316 393994 224368 394000
rect 224144 392142 224264 392170
rect 224144 354550 224172 392142
rect 224224 392080 224276 392086
rect 224224 392022 224276 392028
rect 224236 355502 224264 392022
rect 224224 355496 224276 355502
rect 224224 355438 224276 355444
rect 224132 354544 224184 354550
rect 224132 354486 224184 354492
rect 224040 354476 224092 354482
rect 224040 354418 224092 354424
rect 223948 6452 224000 6458
rect 223948 6394 224000 6400
rect 223856 6384 223908 6390
rect 223856 6326 223908 6332
rect 223764 6316 223816 6322
rect 223764 6258 223816 6264
rect 223488 5228 223540 5234
rect 223488 5170 223540 5176
rect 224328 4146 224356 393994
rect 224408 393916 224460 393922
rect 224408 393858 224460 393864
rect 224420 5370 224448 393858
rect 224696 392086 224724 400044
rect 224788 394058 224816 400044
rect 224880 394126 224908 400044
rect 224972 397905 225000 400044
rect 225064 398138 225092 400044
rect 225052 398132 225104 398138
rect 225052 398074 225104 398080
rect 224958 397896 225014 397905
rect 224958 397831 225014 397840
rect 225156 397633 225184 400044
rect 225142 397624 225198 397633
rect 224960 397588 225012 397594
rect 225142 397559 225198 397568
rect 224960 397530 225012 397536
rect 224868 394120 224920 394126
rect 224868 394062 224920 394068
rect 224776 394052 224828 394058
rect 224776 393994 224828 394000
rect 224684 392080 224736 392086
rect 224684 392022 224736 392028
rect 224972 89010 225000 397530
rect 225052 397520 225104 397526
rect 225248 397497 225276 400044
rect 225340 397730 225368 400044
rect 225432 397769 225460 400044
rect 225418 397760 225474 397769
rect 225328 397724 225380 397730
rect 225418 397695 225474 397704
rect 225328 397666 225380 397672
rect 225052 397462 225104 397468
rect 225234 397488 225290 397497
rect 225064 394058 225092 397462
rect 225234 397423 225290 397432
rect 225524 397322 225552 400044
rect 225616 397526 225644 400044
rect 225604 397520 225656 397526
rect 225604 397462 225656 397468
rect 225512 397316 225564 397322
rect 225512 397258 225564 397264
rect 225708 397202 225736 400044
rect 225156 397174 225736 397202
rect 225052 394052 225104 394058
rect 225052 393994 225104 394000
rect 224960 89004 225012 89010
rect 224960 88946 225012 88952
rect 225156 6526 225184 397174
rect 225800 397066 225828 400044
rect 225340 397038 225828 397066
rect 225236 392012 225288 392018
rect 225236 391954 225288 391960
rect 225144 6520 225196 6526
rect 225144 6462 225196 6468
rect 224408 5364 224460 5370
rect 224408 5306 224460 5312
rect 224316 4140 224368 4146
rect 224316 4082 224368 4088
rect 222844 3868 222896 3874
rect 222844 3810 222896 3816
rect 223948 3528 224000 3534
rect 222304 3454 222792 3482
rect 225248 3482 225276 391954
rect 225340 16182 225368 397038
rect 225892 396930 225920 400044
rect 225432 396902 225920 396930
rect 225432 354618 225460 396902
rect 225984 396794 226012 400044
rect 226076 397390 226104 400044
rect 226064 397384 226116 397390
rect 226064 397326 226116 397332
rect 225524 396766 226012 396794
rect 225420 354612 225472 354618
rect 225420 354554 225472 354560
rect 225328 16176 225380 16182
rect 225328 16118 225380 16124
rect 225524 5438 225552 396766
rect 225788 396704 225840 396710
rect 225788 396646 225840 396652
rect 225604 394664 225656 394670
rect 225604 394606 225656 394612
rect 225512 5432 225564 5438
rect 225512 5374 225564 5380
rect 225616 3942 225644 394606
rect 225800 4826 225828 396646
rect 226168 393314 226196 400044
rect 226260 396710 226288 400044
rect 226352 397497 226380 400044
rect 226444 398410 226472 400044
rect 226432 398404 226484 398410
rect 226432 398346 226484 398352
rect 226536 397633 226564 400044
rect 226522 397624 226578 397633
rect 226522 397559 226578 397568
rect 226432 397520 226484 397526
rect 226338 397488 226394 397497
rect 226432 397462 226484 397468
rect 226338 397423 226394 397432
rect 226248 396704 226300 396710
rect 226248 396646 226300 396652
rect 225892 393286 226196 393314
rect 225892 392766 225920 393286
rect 225880 392760 225932 392766
rect 225880 392702 225932 392708
rect 225788 4820 225840 4826
rect 225788 4762 225840 4768
rect 225604 3936 225656 3942
rect 225604 3878 225656 3884
rect 226444 3534 226472 397462
rect 226628 397458 226656 400044
rect 226616 397452 226668 397458
rect 226616 397394 226668 397400
rect 226720 396778 226748 400044
rect 226708 396772 226760 396778
rect 226708 396714 226760 396720
rect 226812 396658 226840 400044
rect 226628 396630 226840 396658
rect 226524 395344 226576 395350
rect 226524 395286 226576 395292
rect 226536 4010 226564 395286
rect 226524 4004 226576 4010
rect 226524 3946 226576 3952
rect 226628 3738 226656 396630
rect 226708 396568 226760 396574
rect 226708 396510 226760 396516
rect 226720 351218 226748 396510
rect 226800 396500 226852 396506
rect 226800 396442 226852 396448
rect 226812 351966 226840 396442
rect 226904 395350 226932 400044
rect 226892 395344 226944 395350
rect 226892 395286 226944 395292
rect 226996 393314 227024 400044
rect 227088 394670 227116 400044
rect 227180 397594 227208 400044
rect 227168 397588 227220 397594
rect 227168 397530 227220 397536
rect 227168 396772 227220 396778
rect 227168 396714 227220 396720
rect 227076 394664 227128 394670
rect 227076 394606 227128 394612
rect 226904 393286 227024 393314
rect 226800 351960 226852 351966
rect 226800 351902 226852 351908
rect 226708 351212 226760 351218
rect 226708 351154 226760 351160
rect 226904 3806 226932 393286
rect 227180 4078 227208 396714
rect 227272 396574 227300 400044
rect 227260 396568 227312 396574
rect 227260 396510 227312 396516
rect 227364 396370 227392 400044
rect 227456 397798 227484 400044
rect 227444 397792 227496 397798
rect 227444 397734 227496 397740
rect 227548 396506 227576 400044
rect 227640 397662 227668 400044
rect 227628 397656 227680 397662
rect 227628 397598 227680 397604
rect 227732 397526 227760 400044
rect 227720 397520 227772 397526
rect 227720 397462 227772 397468
rect 227824 397186 227852 400044
rect 227812 397180 227864 397186
rect 227812 397122 227864 397128
rect 227812 397044 227864 397050
rect 227812 396986 227864 396992
rect 227536 396500 227588 396506
rect 227536 396442 227588 396448
rect 227352 396364 227404 396370
rect 227352 396306 227404 396312
rect 227168 4072 227220 4078
rect 227168 4014 227220 4020
rect 226892 3800 226944 3806
rect 226892 3742 226944 3748
rect 226616 3732 226668 3738
rect 226616 3674 226668 3680
rect 227824 3670 227852 396986
rect 227916 396710 227944 400044
rect 227904 396704 227956 396710
rect 227904 396646 227956 396652
rect 227904 396568 227956 396574
rect 227904 396510 227956 396516
rect 227916 4146 227944 396510
rect 227904 4140 227956 4146
rect 227904 4082 227956 4088
rect 227812 3664 227864 3670
rect 227812 3606 227864 3612
rect 228008 3534 228036 400044
rect 228100 396914 228128 400044
rect 228088 396908 228140 396914
rect 228088 396850 228140 396856
rect 228192 396794 228220 400044
rect 228284 397730 228312 400044
rect 228272 397724 228324 397730
rect 228272 397666 228324 397672
rect 228100 396766 228220 396794
rect 228100 396574 228128 396766
rect 228180 396704 228232 396710
rect 228180 396646 228232 396652
rect 228272 396704 228324 396710
rect 228272 396646 228324 396652
rect 228088 396568 228140 396574
rect 228088 396510 228140 396516
rect 228088 396432 228140 396438
rect 228088 396374 228140 396380
rect 228100 3738 228128 396374
rect 228088 3732 228140 3738
rect 228088 3674 228140 3680
rect 223948 3470 224000 3476
rect 222764 480 222792 3454
rect 223960 480 223988 3470
rect 225156 3454 225276 3482
rect 226432 3528 226484 3534
rect 226432 3470 226484 3476
rect 227536 3528 227588 3534
rect 227536 3470 227588 3476
rect 227996 3528 228048 3534
rect 227996 3470 228048 3476
rect 225156 480 225184 3454
rect 226340 3188 226392 3194
rect 226340 3130 226392 3136
rect 226352 480 226380 3130
rect 227548 480 227576 3470
rect 228192 3194 228220 396646
rect 228284 177410 228312 396646
rect 228376 394738 228404 400044
rect 228468 398546 228496 400044
rect 228456 398540 228508 398546
rect 228456 398482 228508 398488
rect 228364 394732 228416 394738
rect 228364 394674 228416 394680
rect 228560 393314 228588 400044
rect 228652 396438 228680 400044
rect 228744 397050 228772 400044
rect 228732 397044 228784 397050
rect 228732 396986 228784 396992
rect 228732 396908 228784 396914
rect 228732 396850 228784 396856
rect 228640 396432 228692 396438
rect 228640 396374 228692 396380
rect 228376 393286 228588 393314
rect 228272 177404 228324 177410
rect 228272 177346 228324 177352
rect 228376 177342 228404 393286
rect 228364 177336 228416 177342
rect 228364 177278 228416 177284
rect 228180 3188 228232 3194
rect 228180 3130 228232 3136
rect 228744 480 228772 396850
rect 228836 396710 228864 400044
rect 228928 397497 228956 400044
rect 229020 397633 229048 400044
rect 229006 397624 229062 397633
rect 229006 397559 229062 397568
rect 228914 397488 228970 397497
rect 228914 397423 228970 397432
rect 229008 397180 229060 397186
rect 229008 397122 229060 397128
rect 228824 396704 228876 396710
rect 228824 396646 228876 396652
rect 229020 392018 229048 397122
rect 229112 396438 229140 400044
rect 229204 398177 229232 400044
rect 229296 398834 229324 400044
rect 229388 398993 229416 400044
rect 229374 398984 229430 398993
rect 229374 398919 229430 398928
rect 229296 398806 229416 398834
rect 229284 398676 229336 398682
rect 229284 398618 229336 398624
rect 229190 398168 229246 398177
rect 229190 398103 229246 398112
rect 229296 396794 229324 398618
rect 229388 396846 229416 398806
rect 229204 396766 229324 396794
rect 229376 396840 229428 396846
rect 229376 396782 229428 396788
rect 229100 396432 229152 396438
rect 229100 396374 229152 396380
rect 229008 392012 229060 392018
rect 229008 391954 229060 391960
rect 229204 3466 229232 396766
rect 229480 396658 229508 400044
rect 229572 396778 229600 400044
rect 229560 396772 229612 396778
rect 229560 396714 229612 396720
rect 229664 396658 229692 400044
rect 229756 398342 229784 400044
rect 229744 398336 229796 398342
rect 229744 398278 229796 398284
rect 229742 398168 229798 398177
rect 229742 398103 229798 398112
rect 229756 396982 229784 398103
rect 229744 396976 229796 396982
rect 229744 396918 229796 396924
rect 229296 396630 229508 396658
rect 229572 396630 229692 396658
rect 229192 3460 229244 3466
rect 229192 3402 229244 3408
rect 229296 3398 229324 396630
rect 229376 396568 229428 396574
rect 229376 396510 229428 396516
rect 229388 4894 229416 396510
rect 229468 396500 229520 396506
rect 229468 396442 229520 396448
rect 229376 4888 229428 4894
rect 229376 4830 229428 4836
rect 229480 4826 229508 396442
rect 229572 46238 229600 396630
rect 229652 396432 229704 396438
rect 229652 396374 229704 396380
rect 229664 354006 229692 396374
rect 229848 393314 229876 400044
rect 229940 396506 229968 400044
rect 230032 398682 230060 400044
rect 230020 398676 230072 398682
rect 230020 398618 230072 398624
rect 230020 398540 230072 398546
rect 230020 398482 230072 398488
rect 229928 396500 229980 396506
rect 229928 396442 229980 396448
rect 229756 393286 229876 393314
rect 229756 391270 229784 393286
rect 229744 391264 229796 391270
rect 229744 391206 229796 391212
rect 230032 389978 230060 398482
rect 230124 397633 230152 400044
rect 230216 397905 230244 400044
rect 230202 397896 230258 397905
rect 230202 397831 230258 397840
rect 230110 397624 230166 397633
rect 230110 397559 230166 397568
rect 230308 397497 230336 400044
rect 230400 397769 230428 400044
rect 230492 397882 230520 400044
rect 230584 398274 230612 400044
rect 230572 398268 230624 398274
rect 230572 398210 230624 398216
rect 230492 397854 230612 397882
rect 230386 397760 230442 397769
rect 230386 397695 230442 397704
rect 230480 397724 230532 397730
rect 230480 397666 230532 397672
rect 230294 397488 230350 397497
rect 230294 397423 230350 397432
rect 230112 396840 230164 396846
rect 230112 396782 230164 396788
rect 230020 389972 230072 389978
rect 230020 389914 230072 389920
rect 229652 354000 229704 354006
rect 229652 353942 229704 353948
rect 229560 46232 229612 46238
rect 229560 46174 229612 46180
rect 229468 4820 229520 4826
rect 229468 4762 229520 4768
rect 229836 4140 229888 4146
rect 229836 4082 229888 4088
rect 229284 3392 229336 3398
rect 229284 3334 229336 3340
rect 229848 480 229876 4082
rect 230124 3602 230152 396782
rect 230112 3596 230164 3602
rect 230112 3538 230164 3544
rect 230492 3482 230520 397666
rect 230584 396914 230612 397854
rect 230572 396908 230624 396914
rect 230572 396850 230624 396856
rect 230676 396794 230704 400044
rect 230584 396766 230704 396794
rect 230584 4214 230612 396766
rect 230768 396658 230796 400044
rect 230860 398818 230888 400044
rect 230848 398812 230900 398818
rect 230848 398754 230900 398760
rect 230676 396630 230796 396658
rect 230676 5234 230704 396630
rect 230952 396522 230980 400044
rect 231044 396778 231072 400044
rect 231032 396772 231084 396778
rect 231032 396714 231084 396720
rect 231136 396658 231164 400044
rect 230768 396494 230980 396522
rect 231044 396630 231164 396658
rect 230768 12238 230796 396494
rect 230848 396432 230900 396438
rect 230848 396374 230900 396380
rect 230860 19174 230888 396374
rect 230940 396364 230992 396370
rect 230940 396306 230992 396312
rect 230952 352918 230980 396306
rect 231044 392970 231072 396630
rect 231228 396438 231256 400044
rect 231216 396432 231268 396438
rect 231216 396374 231268 396380
rect 231320 395826 231348 400044
rect 231412 396370 231440 400044
rect 231504 397526 231532 400044
rect 231596 397769 231624 400044
rect 231582 397760 231638 397769
rect 231582 397695 231638 397704
rect 231492 397520 231544 397526
rect 231688 397497 231716 400044
rect 231780 397633 231808 400044
rect 231766 397624 231822 397633
rect 231766 397559 231822 397568
rect 231492 397462 231544 397468
rect 231674 397488 231730 397497
rect 231674 397423 231730 397432
rect 231872 397050 231900 400044
rect 231964 397730 231992 400044
rect 231952 397724 232004 397730
rect 231952 397666 232004 397672
rect 231860 397044 231912 397050
rect 231860 396986 231912 396992
rect 231584 396908 231636 396914
rect 231584 396850 231636 396856
rect 231860 396908 231912 396914
rect 231860 396850 231912 396856
rect 231492 396772 231544 396778
rect 231492 396714 231544 396720
rect 231400 396364 231452 396370
rect 231400 396306 231452 396312
rect 231504 395894 231532 396714
rect 231596 395962 231624 396850
rect 231584 395956 231636 395962
rect 231584 395898 231636 395904
rect 231492 395888 231544 395894
rect 231492 395830 231544 395836
rect 231308 395820 231360 395826
rect 231308 395762 231360 395768
rect 231124 394732 231176 394738
rect 231124 394674 231176 394680
rect 231032 392964 231084 392970
rect 231032 392906 231084 392912
rect 230940 352912 230992 352918
rect 230940 352854 230992 352860
rect 230848 19168 230900 19174
rect 230848 19110 230900 19116
rect 230756 12232 230808 12238
rect 230756 12174 230808 12180
rect 230664 5228 230716 5234
rect 230664 5170 230716 5176
rect 230572 4208 230624 4214
rect 230572 4150 230624 4156
rect 231136 3534 231164 394674
rect 231872 6526 231900 396850
rect 231952 396840 232004 396846
rect 231952 396782 232004 396788
rect 231964 18970 231992 396782
rect 232056 19038 232084 400044
rect 232148 396658 232176 400044
rect 232240 396778 232268 400044
rect 232332 396846 232360 400044
rect 232320 396840 232372 396846
rect 232320 396782 232372 396788
rect 232228 396772 232280 396778
rect 232228 396714 232280 396720
rect 232148 396630 232360 396658
rect 232228 396568 232280 396574
rect 232134 396536 232190 396545
rect 232228 396510 232280 396516
rect 232134 396471 232190 396480
rect 232148 20262 232176 396471
rect 232240 25906 232268 396510
rect 232332 25974 232360 396630
rect 232424 396574 232452 400044
rect 232516 396914 232544 400044
rect 232504 396908 232556 396914
rect 232504 396850 232556 396856
rect 232608 396817 232636 400044
rect 232594 396808 232650 396817
rect 232700 396778 232728 400044
rect 232594 396743 232650 396752
rect 232688 396772 232740 396778
rect 232688 396714 232740 396720
rect 232792 396658 232820 400044
rect 232884 397633 232912 400044
rect 232976 397905 233004 400044
rect 232962 397896 233018 397905
rect 232962 397831 233018 397840
rect 232870 397624 232926 397633
rect 232870 397559 232926 397568
rect 233068 397497 233096 400044
rect 233160 397769 233188 400044
rect 233146 397760 233202 397769
rect 233146 397695 233202 397704
rect 233054 397488 233110 397497
rect 233054 397423 233110 397432
rect 232872 397044 232924 397050
rect 232872 396986 232924 396992
rect 232516 396630 232820 396658
rect 232412 396568 232464 396574
rect 232412 396510 232464 396516
rect 232412 396432 232464 396438
rect 232412 396374 232464 396380
rect 232424 87786 232452 396374
rect 232516 355570 232544 396630
rect 232596 396568 232648 396574
rect 232596 396510 232648 396516
rect 232608 355638 232636 396510
rect 232884 395758 232912 396986
rect 233252 396370 233280 400044
rect 233344 398478 233372 400044
rect 233332 398472 233384 398478
rect 233332 398414 233384 398420
rect 233332 396908 233384 396914
rect 233332 396850 233384 396856
rect 233344 396522 233372 396850
rect 233436 396658 233464 400044
rect 233528 396794 233556 400044
rect 233620 398546 233648 400044
rect 233608 398540 233660 398546
rect 233608 398482 233660 398488
rect 233712 396914 233740 400044
rect 233700 396908 233752 396914
rect 233700 396850 233752 396856
rect 233528 396766 233740 396794
rect 233436 396630 233648 396658
rect 233516 396568 233568 396574
rect 233344 396494 233464 396522
rect 233516 396510 233568 396516
rect 233332 396432 233384 396438
rect 233332 396374 233384 396380
rect 233240 396364 233292 396370
rect 233240 396306 233292 396312
rect 233240 396228 233292 396234
rect 233240 396170 233292 396176
rect 232872 395752 232924 395758
rect 232872 395694 232924 395700
rect 232596 355632 232648 355638
rect 232596 355574 232648 355580
rect 232504 355564 232556 355570
rect 232504 355506 232556 355512
rect 232504 177404 232556 177410
rect 232504 177346 232556 177352
rect 232412 87780 232464 87786
rect 232412 87722 232464 87728
rect 232320 25968 232372 25974
rect 232320 25910 232372 25916
rect 232228 25900 232280 25906
rect 232228 25842 232280 25848
rect 232136 20256 232188 20262
rect 232136 20198 232188 20204
rect 232044 19032 232096 19038
rect 232044 18974 232096 18980
rect 231952 18964 232004 18970
rect 231952 18906 232004 18912
rect 231860 6520 231912 6526
rect 231860 6462 231912 6468
rect 231124 3528 231176 3534
rect 230492 3454 231072 3482
rect 231124 3470 231176 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 231044 480 231072 3454
rect 232240 480 232268 3470
rect 232516 3126 232544 177346
rect 233252 7886 233280 396170
rect 233344 7954 233372 396374
rect 233436 391474 233464 396494
rect 233424 391468 233476 391474
rect 233424 391410 233476 391416
rect 233424 389972 233476 389978
rect 233424 389914 233476 389920
rect 233332 7948 233384 7954
rect 233332 7890 233384 7896
rect 233240 7880 233292 7886
rect 233240 7822 233292 7828
rect 232504 3120 232556 3126
rect 232504 3062 232556 3068
rect 233436 480 233464 389914
rect 233528 18902 233556 396510
rect 233620 20194 233648 396630
rect 233712 83638 233740 396766
rect 233804 351354 233832 400044
rect 233896 396438 233924 400044
rect 233988 396574 234016 400044
rect 234080 397662 234108 400044
rect 234068 397656 234120 397662
rect 234068 397598 234120 397604
rect 234068 397520 234120 397526
rect 234068 397462 234120 397468
rect 233976 396568 234028 396574
rect 233976 396510 234028 396516
rect 233884 396432 233936 396438
rect 233884 396374 233936 396380
rect 233976 396364 234028 396370
rect 233976 396306 234028 396312
rect 233884 396296 233936 396302
rect 233884 396238 233936 396244
rect 233792 351348 233844 351354
rect 233792 351290 233844 351296
rect 233700 83632 233752 83638
rect 233700 83574 233752 83580
rect 233608 20188 233660 20194
rect 233608 20130 233660 20136
rect 233896 19106 233924 396238
rect 233988 390046 234016 396306
rect 234080 396302 234108 397462
rect 234068 396296 234120 396302
rect 234068 396238 234120 396244
rect 234172 396234 234200 400044
rect 234264 397497 234292 400044
rect 234356 397633 234384 400044
rect 234448 397769 234476 400044
rect 234434 397760 234490 397769
rect 234434 397695 234490 397704
rect 234342 397624 234398 397633
rect 234342 397559 234398 397568
rect 234344 397520 234396 397526
rect 234250 397488 234306 397497
rect 234540 397474 234568 400044
rect 234344 397462 234396 397468
rect 234250 397423 234306 397432
rect 234160 396228 234212 396234
rect 234160 396170 234212 396176
rect 234356 394534 234384 397462
rect 234448 397446 234568 397474
rect 234448 396545 234476 397446
rect 234632 397066 234660 400044
rect 234724 399945 234752 400044
rect 234710 399936 234766 399945
rect 234710 399871 234766 399880
rect 234816 397066 234844 400044
rect 234540 397038 234660 397066
rect 234724 397038 234844 397066
rect 234908 397050 234936 400044
rect 234896 397044 234948 397050
rect 234540 396574 234568 397038
rect 234620 396908 234672 396914
rect 234620 396850 234672 396856
rect 234528 396568 234580 396574
rect 234434 396536 234490 396545
rect 234528 396510 234580 396516
rect 234434 396471 234490 396480
rect 234344 394528 234396 394534
rect 234344 394470 234396 394476
rect 233976 390040 234028 390046
rect 233976 389982 234028 389988
rect 233884 19100 233936 19106
rect 233884 19042 233936 19048
rect 233516 18896 233568 18902
rect 233516 18838 233568 18844
rect 234632 7818 234660 396850
rect 234724 396658 234752 397038
rect 234896 396986 234948 396992
rect 235000 396914 235028 400044
rect 234988 396908 235040 396914
rect 234988 396850 235040 396856
rect 234988 396772 235040 396778
rect 234988 396714 235040 396720
rect 234724 396630 234936 396658
rect 234804 396500 234856 396506
rect 234804 396442 234856 396448
rect 234816 9314 234844 396442
rect 234908 20126 234936 396630
rect 235000 25770 235028 396714
rect 235092 396658 235120 400044
rect 235184 396778 235212 400044
rect 235276 396778 235304 400044
rect 235172 396772 235224 396778
rect 235172 396714 235224 396720
rect 235264 396772 235316 396778
rect 235264 396714 235316 396720
rect 235368 396658 235396 400044
rect 235460 397186 235488 400044
rect 235448 397180 235500 397186
rect 235448 397122 235500 397128
rect 235448 397044 235500 397050
rect 235448 396986 235500 396992
rect 235092 396630 235212 396658
rect 235080 396568 235132 396574
rect 235080 396510 235132 396516
rect 235092 25838 235120 396510
rect 235184 352850 235212 396630
rect 235276 396630 235396 396658
rect 235172 352844 235224 352850
rect 235172 352786 235224 352792
rect 235276 352782 235304 396630
rect 235460 393314 235488 396986
rect 235552 396506 235580 400044
rect 235644 397361 235672 400044
rect 235736 397633 235764 400044
rect 235722 397624 235778 397633
rect 235722 397559 235778 397568
rect 235828 397497 235856 400044
rect 235920 397769 235948 400044
rect 235906 397760 235962 397769
rect 235906 397695 235962 397704
rect 235814 397488 235870 397497
rect 235814 397423 235870 397432
rect 235630 397352 235686 397361
rect 235630 397287 235686 397296
rect 235632 397180 235684 397186
rect 235632 397122 235684 397128
rect 235540 396500 235592 396506
rect 235540 396442 235592 396448
rect 235644 394466 235672 397122
rect 235908 396772 235960 396778
rect 235908 396714 235960 396720
rect 235632 394460 235684 394466
rect 235632 394402 235684 394408
rect 235368 393286 235488 393314
rect 235368 389978 235396 393286
rect 235356 389972 235408 389978
rect 235356 389914 235408 389920
rect 235264 352776 235316 352782
rect 235264 352718 235316 352724
rect 235172 177336 235224 177342
rect 235172 177278 235224 177284
rect 235080 25832 235132 25838
rect 235080 25774 235132 25780
rect 234988 25764 235040 25770
rect 234988 25706 235040 25712
rect 234896 20120 234948 20126
rect 234896 20062 234948 20068
rect 234804 9308 234856 9314
rect 234804 9250 234856 9256
rect 234620 7812 234672 7818
rect 234620 7754 234672 7760
rect 235184 6914 235212 177278
rect 235920 7750 235948 396714
rect 236012 396522 236040 400044
rect 236104 398954 236132 400044
rect 236092 398948 236144 398954
rect 236092 398890 236144 398896
rect 236196 396658 236224 400044
rect 236288 396778 236316 400044
rect 236380 397866 236408 400044
rect 236368 397860 236420 397866
rect 236368 397802 236420 397808
rect 236276 396772 236328 396778
rect 236276 396714 236328 396720
rect 236368 396704 236420 396710
rect 236196 396630 236316 396658
rect 236368 396646 236420 396652
rect 236012 396494 236224 396522
rect 236092 396432 236144 396438
rect 236092 396374 236144 396380
rect 236000 396364 236052 396370
rect 236000 396306 236052 396312
rect 236012 9178 236040 396306
rect 236104 9246 236132 396374
rect 236196 12170 236224 396494
rect 236288 20058 236316 396630
rect 236380 21690 236408 396646
rect 236472 21758 236500 400044
rect 236564 80714 236592 400044
rect 236656 396438 236684 400044
rect 236748 396710 236776 400044
rect 236736 396704 236788 396710
rect 236736 396646 236788 396652
rect 236644 396432 236696 396438
rect 236644 396374 236696 396380
rect 236840 394330 236868 400044
rect 236932 396370 236960 400044
rect 237024 396914 237052 400044
rect 237116 397769 237144 400044
rect 237102 397760 237158 397769
rect 237102 397695 237158 397704
rect 237208 397497 237236 400044
rect 237300 397633 237328 400044
rect 237286 397624 237342 397633
rect 237286 397559 237342 397568
rect 237194 397488 237250 397497
rect 237194 397423 237250 397432
rect 237392 396982 237420 400044
rect 237380 396976 237432 396982
rect 237380 396918 237432 396924
rect 237012 396908 237064 396914
rect 237012 396850 237064 396856
rect 237012 396772 237064 396778
rect 237012 396714 237064 396720
rect 237380 396772 237432 396778
rect 237380 396714 237432 396720
rect 236920 396364 236972 396370
rect 236920 396306 236972 396312
rect 237024 394398 237052 396714
rect 237012 394392 237064 394398
rect 237012 394334 237064 394340
rect 236828 394324 236880 394330
rect 236828 394266 236880 394272
rect 236552 80708 236604 80714
rect 236552 80650 236604 80656
rect 236460 21752 236512 21758
rect 236460 21694 236512 21700
rect 236368 21684 236420 21690
rect 236368 21626 236420 21632
rect 236276 20052 236328 20058
rect 236276 19994 236328 20000
rect 236184 12164 236236 12170
rect 236184 12106 236236 12112
rect 236092 9240 236144 9246
rect 236092 9182 236144 9188
rect 236000 9172 236052 9178
rect 236000 9114 236052 9120
rect 237392 9042 237420 396714
rect 237484 9110 237512 400044
rect 237576 396370 237604 400044
rect 237668 396658 237696 400044
rect 237760 396778 237788 400044
rect 237748 396772 237800 396778
rect 237748 396714 237800 396720
rect 237668 396630 237788 396658
rect 237656 396568 237708 396574
rect 237656 396510 237708 396516
rect 237564 396364 237616 396370
rect 237564 396306 237616 396312
rect 237668 396250 237696 396510
rect 237576 396222 237696 396250
rect 237472 9104 237524 9110
rect 237472 9046 237524 9052
rect 237380 9036 237432 9042
rect 237380 8978 237432 8984
rect 237576 8974 237604 396222
rect 237656 396160 237708 396166
rect 237656 396102 237708 396108
rect 237668 10674 237696 396102
rect 237760 13462 237788 396630
rect 237852 396522 237880 400044
rect 237944 396658 237972 400044
rect 238036 396778 238064 400044
rect 238024 396772 238076 396778
rect 238024 396714 238076 396720
rect 238128 396658 238156 400044
rect 238220 398002 238248 400044
rect 238208 397996 238260 398002
rect 238208 397938 238260 397944
rect 237944 396630 238064 396658
rect 238128 396630 238248 396658
rect 237852 396506 237972 396522
rect 237852 396500 237984 396506
rect 237852 396494 237932 396500
rect 237932 396442 237984 396448
rect 237840 396432 237892 396438
rect 237840 396374 237892 396380
rect 237852 21554 237880 396374
rect 237932 396364 237984 396370
rect 237932 396306 237984 396312
rect 237944 21622 237972 396306
rect 238036 84862 238064 396630
rect 238116 396500 238168 396506
rect 238116 396442 238168 396448
rect 238128 354346 238156 396442
rect 238220 396438 238248 396630
rect 238208 396432 238260 396438
rect 238208 396374 238260 396380
rect 238312 396166 238340 400044
rect 238404 397497 238432 400044
rect 238496 397633 238524 400044
rect 238588 397769 238616 400044
rect 238574 397760 238630 397769
rect 238574 397695 238630 397704
rect 238482 397624 238538 397633
rect 238482 397559 238538 397568
rect 238390 397488 238446 397497
rect 238390 397423 238446 397432
rect 238680 397225 238708 400044
rect 238772 397526 238800 400044
rect 238760 397520 238812 397526
rect 238760 397462 238812 397468
rect 238666 397216 238722 397225
rect 238666 397151 238722 397160
rect 238760 397180 238812 397186
rect 238760 397122 238812 397128
rect 238392 396976 238444 396982
rect 238392 396918 238444 396924
rect 238300 396160 238352 396166
rect 238300 396102 238352 396108
rect 238404 394262 238432 396918
rect 238392 394256 238444 394262
rect 238392 394198 238444 394204
rect 238116 354340 238168 354346
rect 238116 354282 238168 354288
rect 238024 84856 238076 84862
rect 238024 84798 238076 84804
rect 237932 21616 237984 21622
rect 237932 21558 237984 21564
rect 237840 21548 237892 21554
rect 237840 21490 237892 21496
rect 237748 13456 237800 13462
rect 237748 13398 237800 13404
rect 237656 10668 237708 10674
rect 237656 10610 237708 10616
rect 238772 10538 238800 397122
rect 238864 397050 238892 400044
rect 238852 397044 238904 397050
rect 238852 396986 238904 396992
rect 238956 396982 238984 400044
rect 238944 396976 238996 396982
rect 238944 396918 238996 396924
rect 238850 396808 238906 396817
rect 239048 396794 239076 400044
rect 239140 396817 239168 400044
rect 238850 396743 238906 396752
rect 238956 396766 239076 396794
rect 239126 396808 239182 396817
rect 238864 10606 238892 396743
rect 238956 14822 238984 396766
rect 239126 396743 239182 396752
rect 239128 396704 239180 396710
rect 239128 396646 239180 396652
rect 239036 396568 239088 396574
rect 239036 396510 239088 396516
rect 239048 16318 239076 396510
rect 239140 21418 239168 396646
rect 239232 21486 239260 400044
rect 239324 398002 239352 400044
rect 239312 397996 239364 398002
rect 239312 397938 239364 397944
rect 239312 397860 239364 397866
rect 239312 397802 239364 397808
rect 239324 397594 239352 397802
rect 239312 397588 239364 397594
rect 239312 397530 239364 397536
rect 239416 397186 239444 400044
rect 239404 397180 239456 397186
rect 239404 397122 239456 397128
rect 239404 397044 239456 397050
rect 239404 396986 239456 396992
rect 239312 396976 239364 396982
rect 239312 396918 239364 396924
rect 239324 352714 239352 396918
rect 239416 391406 239444 396986
rect 239508 396710 239536 400044
rect 239496 396704 239548 396710
rect 239496 396646 239548 396652
rect 239600 396574 239628 400044
rect 239692 397497 239720 400044
rect 239784 397633 239812 400044
rect 239876 398614 239904 400044
rect 239864 398608 239916 398614
rect 239864 398550 239916 398556
rect 239864 398472 239916 398478
rect 239864 398414 239916 398420
rect 239770 397624 239826 397633
rect 239770 397559 239826 397568
rect 239678 397488 239734 397497
rect 239678 397423 239734 397432
rect 239588 396568 239640 396574
rect 239588 396510 239640 396516
rect 239876 393314 239904 398414
rect 239968 397497 239996 400044
rect 240060 397769 240088 400044
rect 240046 397760 240102 397769
rect 240046 397695 240102 397704
rect 240048 397588 240100 397594
rect 240048 397530 240100 397536
rect 239954 397488 240010 397497
rect 239954 397423 240010 397432
rect 240060 395690 240088 397530
rect 240152 396794 240180 400044
rect 240244 399945 240272 400044
rect 240230 399936 240286 399945
rect 240230 399871 240286 399880
rect 240152 396766 240272 396794
rect 240336 396778 240364 400044
rect 240428 398478 240456 400044
rect 240416 398472 240468 398478
rect 240416 398414 240468 398420
rect 240140 396500 240192 396506
rect 240140 396442 240192 396448
rect 240048 395684 240100 395690
rect 240048 395626 240100 395632
rect 239600 393286 239904 393314
rect 239600 392902 239628 393286
rect 239588 392896 239640 392902
rect 239588 392838 239640 392844
rect 239404 391400 239456 391406
rect 239404 391342 239456 391348
rect 239312 352708 239364 352714
rect 239312 352650 239364 352656
rect 239220 21480 239272 21486
rect 239220 21422 239272 21428
rect 239128 21412 239180 21418
rect 239128 21354 239180 21360
rect 239036 16312 239088 16318
rect 239036 16254 239088 16260
rect 238944 14816 238996 14822
rect 238944 14758 238996 14764
rect 238852 10600 238904 10606
rect 238852 10542 238904 10548
rect 238760 10532 238812 10538
rect 238760 10474 238812 10480
rect 237564 8968 237616 8974
rect 237564 8910 237616 8916
rect 235908 7744 235960 7750
rect 235908 7686 235960 7692
rect 234632 6886 235212 6914
rect 234632 480 234660 6886
rect 240152 6458 240180 396442
rect 240244 394126 240272 396766
rect 240324 396772 240376 396778
rect 240324 396714 240376 396720
rect 240520 396658 240548 400044
rect 240612 396778 240640 400044
rect 240600 396772 240652 396778
rect 240600 396714 240652 396720
rect 240704 396658 240732 400044
rect 240796 396982 240824 400044
rect 240784 396976 240836 396982
rect 240784 396918 240836 396924
rect 240784 396772 240836 396778
rect 240784 396714 240836 396720
rect 240428 396630 240548 396658
rect 240612 396630 240732 396658
rect 240428 396506 240456 396630
rect 240416 396500 240468 396506
rect 240416 396442 240468 396448
rect 240508 396500 240560 396506
rect 240508 396442 240560 396448
rect 240324 396432 240376 396438
rect 240324 396374 240376 396380
rect 240232 394120 240284 394126
rect 240232 394062 240284 394068
rect 240336 10402 240364 396374
rect 240416 396364 240468 396370
rect 240416 396306 240468 396312
rect 240428 17610 240456 396306
rect 240520 18834 240548 396442
rect 240612 25702 240640 396630
rect 240692 396568 240744 396574
rect 240692 396510 240744 396516
rect 240704 86358 240732 396510
rect 240796 178702 240824 396714
rect 240888 354278 240916 400044
rect 240980 397526 241008 400044
rect 240968 397520 241020 397526
rect 240968 397462 241020 397468
rect 241072 396438 241100 400044
rect 241164 396506 241192 400044
rect 241152 396500 241204 396506
rect 241152 396442 241204 396448
rect 241060 396432 241112 396438
rect 241060 396374 241112 396380
rect 241256 396370 241284 400044
rect 241348 397497 241376 400044
rect 241334 397488 241390 397497
rect 241334 397423 241390 397432
rect 241440 397089 241468 400044
rect 241532 398342 241560 400044
rect 241520 398336 241572 398342
rect 241520 398278 241572 398284
rect 241426 397080 241482 397089
rect 241426 397015 241482 397024
rect 241428 396976 241480 396982
rect 241428 396918 241480 396924
rect 241244 396364 241296 396370
rect 241244 396306 241296 396312
rect 240876 354272 240928 354278
rect 240876 354214 240928 354220
rect 240784 178696 240836 178702
rect 240784 178638 240836 178644
rect 240692 86352 240744 86358
rect 240692 86294 240744 86300
rect 240600 25696 240652 25702
rect 240600 25638 240652 25644
rect 240508 18828 240560 18834
rect 240508 18770 240560 18776
rect 240416 17604 240468 17610
rect 240416 17546 240468 17552
rect 241440 10470 241468 396918
rect 241520 396772 241572 396778
rect 241520 396714 241572 396720
rect 241532 12034 241560 396714
rect 241624 396522 241652 400044
rect 241716 397186 241744 400044
rect 241704 397180 241756 397186
rect 241704 397122 241756 397128
rect 241808 396658 241836 400044
rect 241900 396778 241928 400044
rect 241888 396772 241940 396778
rect 241888 396714 241940 396720
rect 241808 396630 241928 396658
rect 241624 396494 241836 396522
rect 241704 396432 241756 396438
rect 241704 396374 241756 396380
rect 241612 396364 241664 396370
rect 241612 396306 241664 396312
rect 241520 12028 241572 12034
rect 241520 11970 241572 11976
rect 241624 11966 241652 396306
rect 241716 23050 241744 396374
rect 241808 392834 241836 396494
rect 241796 392828 241848 392834
rect 241796 392770 241848 392776
rect 241796 354000 241848 354006
rect 241796 353942 241848 353948
rect 241704 23044 241756 23050
rect 241704 22986 241756 22992
rect 241612 11960 241664 11966
rect 241612 11902 241664 11908
rect 241428 10464 241480 10470
rect 241428 10406 241480 10412
rect 240324 10396 240376 10402
rect 240324 10338 240376 10344
rect 241808 6914 241836 353942
rect 241900 352578 241928 396630
rect 241992 396438 242020 400044
rect 242084 398206 242112 400044
rect 242072 398200 242124 398206
rect 242072 398142 242124 398148
rect 241980 396432 242032 396438
rect 241980 396374 242032 396380
rect 242176 396370 242204 400044
rect 242268 396914 242296 400044
rect 242256 396908 242308 396914
rect 242256 396850 242308 396856
rect 242164 396364 242216 396370
rect 242164 396306 242216 396312
rect 242360 393530 242388 400044
rect 242452 397633 242480 400044
rect 242544 397769 242572 400044
rect 242636 398177 242664 400044
rect 242622 398168 242678 398177
rect 242622 398103 242678 398112
rect 242624 397996 242676 398002
rect 242624 397938 242676 397944
rect 242530 397760 242586 397769
rect 242530 397695 242586 397704
rect 242438 397624 242494 397633
rect 242636 397610 242664 397938
rect 242438 397559 242494 397568
rect 242544 397582 242664 397610
rect 242440 396840 242492 396846
rect 242440 396782 242492 396788
rect 241992 393502 242388 393530
rect 241992 354210 242020 393502
rect 242452 393394 242480 396782
rect 242176 393366 242480 393394
rect 241980 354204 242032 354210
rect 241980 354146 242032 354152
rect 241888 352572 241940 352578
rect 241888 352514 241940 352520
rect 241716 6886 241836 6914
rect 240140 6452 240192 6458
rect 240140 6394 240192 6400
rect 237378 5400 237434 5409
rect 237378 5335 237434 5344
rect 235816 3732 235868 3738
rect 235816 3674 235868 3680
rect 235828 480 235856 3674
rect 237392 3670 237420 5335
rect 239310 3768 239366 3777
rect 239310 3703 239366 3712
rect 237012 3664 237064 3670
rect 237012 3606 237064 3612
rect 237380 3664 237432 3670
rect 237380 3606 237432 3612
rect 237024 480 237052 3606
rect 238116 3120 238168 3126
rect 238116 3062 238168 3068
rect 238128 480 238156 3062
rect 239324 480 239352 3703
rect 240506 3632 240562 3641
rect 240506 3567 240562 3576
rect 240520 480 240548 3567
rect 241716 480 241744 6886
rect 242176 3194 242204 393366
rect 242544 393314 242572 397582
rect 242624 397520 242676 397526
rect 242728 397497 242756 400044
rect 242820 397905 242848 400044
rect 242806 397896 242862 397905
rect 242806 397831 242862 397840
rect 242624 397462 242676 397468
rect 242714 397488 242770 397497
rect 242268 393286 242572 393314
rect 242268 177342 242296 393286
rect 242636 351286 242664 397462
rect 242714 397423 242770 397432
rect 242808 396840 242860 396846
rect 242808 396782 242860 396788
rect 242820 396386 242848 396782
rect 242912 396506 242940 400044
rect 242900 396500 242952 396506
rect 242900 396442 242952 396448
rect 242820 396358 242940 396386
rect 242624 351280 242676 351286
rect 242624 351222 242676 351228
rect 242256 177336 242308 177342
rect 242256 177278 242308 177284
rect 242912 11762 242940 396358
rect 243004 11898 243032 400044
rect 243096 396778 243124 400044
rect 243188 397866 243216 400044
rect 243176 397860 243228 397866
rect 243176 397802 243228 397808
rect 243084 396772 243136 396778
rect 243084 396714 243136 396720
rect 243280 396658 243308 400044
rect 243372 396778 243400 400044
rect 243360 396772 243412 396778
rect 243360 396714 243412 396720
rect 243464 396658 243492 400044
rect 243556 396846 243584 400044
rect 243544 396840 243596 396846
rect 243544 396782 243596 396788
rect 243648 396658 243676 400044
rect 243740 397798 243768 400044
rect 243728 397792 243780 397798
rect 243728 397734 243780 397740
rect 243728 396772 243780 396778
rect 243728 396714 243780 396720
rect 243096 396630 243308 396658
rect 243372 396630 243492 396658
rect 243556 396630 243676 396658
rect 242992 11892 243044 11898
rect 242992 11834 243044 11840
rect 243096 11830 243124 396630
rect 243268 396500 243320 396506
rect 243268 396442 243320 396448
rect 243176 396432 243228 396438
rect 243176 396374 243228 396380
rect 243188 13394 243216 396374
rect 243280 18766 243308 396442
rect 243372 25634 243400 396630
rect 243452 396568 243504 396574
rect 243452 396510 243504 396516
rect 243464 83502 243492 396510
rect 243556 87718 243584 396630
rect 243740 393314 243768 396714
rect 243832 396438 243860 400044
rect 243924 396953 243952 400044
rect 244016 397633 244044 400044
rect 244002 397624 244058 397633
rect 244002 397559 244058 397568
rect 244004 397520 244056 397526
rect 244108 397497 244136 400044
rect 244200 397769 244228 400044
rect 244292 398070 244320 400044
rect 244384 399158 244412 400044
rect 244372 399152 244424 399158
rect 244372 399094 244424 399100
rect 244476 398834 244504 400044
rect 244384 398806 244504 398834
rect 244280 398064 244332 398070
rect 244280 398006 244332 398012
rect 244186 397760 244242 397769
rect 244186 397695 244242 397704
rect 244004 397462 244056 397468
rect 244094 397488 244150 397497
rect 243910 396944 243966 396953
rect 243910 396879 243966 396888
rect 243820 396432 243872 396438
rect 243820 396374 243872 396380
rect 244016 394194 244044 397462
rect 244094 397423 244150 397432
rect 244384 396930 244412 398806
rect 244464 397656 244516 397662
rect 244464 397598 244516 397604
rect 244476 397526 244504 397598
rect 244464 397520 244516 397526
rect 244464 397462 244516 397468
rect 244200 396902 244412 396930
rect 244200 396166 244228 396902
rect 244188 396160 244240 396166
rect 244188 396102 244240 396108
rect 244568 394670 244596 400044
rect 244556 394664 244608 394670
rect 244556 394606 244608 394612
rect 244004 394188 244056 394194
rect 244004 394130 244056 394136
rect 244660 393938 244688 400044
rect 243648 393286 243768 393314
rect 244292 393910 244688 393938
rect 243648 351218 243676 393286
rect 243636 351212 243688 351218
rect 243636 351154 243688 351160
rect 243544 87712 243596 87718
rect 243544 87654 243596 87660
rect 243452 83496 243504 83502
rect 243452 83438 243504 83444
rect 243360 25628 243412 25634
rect 243360 25570 243412 25576
rect 243268 18760 243320 18766
rect 243268 18702 243320 18708
rect 243176 13388 243228 13394
rect 243176 13330 243228 13336
rect 244292 13326 244320 393910
rect 244464 393848 244516 393854
rect 244464 393790 244516 393796
rect 244372 393780 244424 393786
rect 244372 393722 244424 393728
rect 244280 13320 244332 13326
rect 244280 13262 244332 13268
rect 244384 13190 244412 393722
rect 244476 13258 244504 393790
rect 244752 393258 244780 400044
rect 244844 398750 244872 400044
rect 244832 398744 244884 398750
rect 244832 398686 244884 398692
rect 244832 397928 244884 397934
rect 244832 397870 244884 397876
rect 244844 397730 244872 397870
rect 244832 397724 244884 397730
rect 244832 397666 244884 397672
rect 244936 394058 244964 400044
rect 244924 394052 244976 394058
rect 244924 393994 244976 394000
rect 245028 393938 245056 400044
rect 244568 393230 244780 393258
rect 244844 393910 245056 393938
rect 244568 22982 244596 393230
rect 244740 393168 244792 393174
rect 244740 393110 244792 393116
rect 244648 393100 244700 393106
rect 244648 393042 244700 393048
rect 244556 22976 244608 22982
rect 244556 22918 244608 22924
rect 244660 22914 244688 393042
rect 244752 26994 244780 393110
rect 244844 354142 244872 393910
rect 245120 393174 245148 400044
rect 245212 393786 245240 400044
rect 245200 393780 245252 393786
rect 245200 393722 245252 393728
rect 245108 393168 245160 393174
rect 245108 393110 245160 393116
rect 245304 393106 245332 400044
rect 245396 398993 245424 400044
rect 245382 398984 245438 398993
rect 245382 398919 245438 398928
rect 245384 398472 245436 398478
rect 245384 398414 245436 398420
rect 245292 393100 245344 393106
rect 245292 393042 245344 393048
rect 245396 389174 245424 398414
rect 245488 397497 245516 400044
rect 245474 397488 245530 397497
rect 245474 397423 245530 397432
rect 245580 396817 245608 400044
rect 245672 398834 245700 400044
rect 245764 399945 245792 400044
rect 245750 399936 245806 399945
rect 245750 399871 245806 399880
rect 245672 398806 245792 398834
rect 245660 398608 245712 398614
rect 245660 398550 245712 398556
rect 245672 398138 245700 398550
rect 245660 398132 245712 398138
rect 245660 398074 245712 398080
rect 245566 396808 245622 396817
rect 245566 396743 245622 396752
rect 245476 396160 245528 396166
rect 245476 396102 245528 396108
rect 245488 389842 245516 396102
rect 245764 396074 245792 398806
rect 245672 396046 245792 396074
rect 245856 396074 245884 400044
rect 245948 398546 245976 400044
rect 245936 398540 245988 398546
rect 245936 398482 245988 398488
rect 245936 397928 245988 397934
rect 245936 397870 245988 397876
rect 245948 397730 245976 397870
rect 245936 397724 245988 397730
rect 245936 397666 245988 397672
rect 245856 396046 245976 396074
rect 245568 394664 245620 394670
rect 245568 394606 245620 394612
rect 245580 393922 245608 394606
rect 245672 394346 245700 396046
rect 245672 394318 245792 394346
rect 245568 393916 245620 393922
rect 245568 393858 245620 393864
rect 245660 392420 245712 392426
rect 245660 392362 245712 392368
rect 245476 389836 245528 389842
rect 245476 389778 245528 389784
rect 244936 389146 245424 389174
rect 244832 354136 244884 354142
rect 244832 354078 244884 354084
rect 244740 26988 244792 26994
rect 244740 26930 244792 26936
rect 244936 23118 244964 389146
rect 244924 23112 244976 23118
rect 244924 23054 244976 23060
rect 244648 22908 244700 22914
rect 244648 22850 244700 22856
rect 244464 13252 244516 13258
rect 244464 13194 244516 13200
rect 244372 13184 244424 13190
rect 244372 13126 244424 13132
rect 245672 13122 245700 392362
rect 245764 391202 245792 394318
rect 245844 393848 245896 393854
rect 245844 393790 245896 393796
rect 245752 391196 245804 391202
rect 245752 391138 245804 391144
rect 245856 14686 245884 393790
rect 245948 22846 245976 396046
rect 246040 392426 246068 400044
rect 246028 392420 246080 392426
rect 246028 392362 246080 392368
rect 246132 392306 246160 400044
rect 246224 398478 246252 400044
rect 246212 398472 246264 398478
rect 246212 398414 246264 398420
rect 246210 398304 246266 398313
rect 246210 398239 246266 398248
rect 246224 397118 246252 398239
rect 246212 397112 246264 397118
rect 246212 397054 246264 397060
rect 246316 393990 246344 400044
rect 246304 393984 246356 393990
rect 246304 393926 246356 393932
rect 246040 392278 246160 392306
rect 245936 22840 245988 22846
rect 245936 22782 245988 22788
rect 246040 22778 246068 392278
rect 246408 392170 246436 400044
rect 246500 398721 246528 400044
rect 246486 398712 246542 398721
rect 246486 398647 246542 398656
rect 246488 398132 246540 398138
rect 246488 398074 246540 398080
rect 246132 392142 246436 392170
rect 246132 24478 246160 392142
rect 246212 391196 246264 391202
rect 246212 391138 246264 391144
rect 246224 86290 246252 391138
rect 246500 389174 246528 398074
rect 246592 393854 246620 400044
rect 246684 397633 246712 400044
rect 246776 397905 246804 400044
rect 246762 397896 246818 397905
rect 246762 397831 246818 397840
rect 246764 397724 246816 397730
rect 246764 397666 246816 397672
rect 246670 397624 246726 397633
rect 246670 397559 246726 397568
rect 246580 393848 246632 393854
rect 246580 393790 246632 393796
rect 246776 389910 246804 397666
rect 246868 397497 246896 400044
rect 246960 397769 246988 400044
rect 246946 397760 247002 397769
rect 246946 397695 247002 397704
rect 246854 397488 246910 397497
rect 246854 397423 246910 397432
rect 247052 397254 247080 400044
rect 247040 397248 247092 397254
rect 247040 397190 247092 397196
rect 247038 397080 247094 397089
rect 247038 397015 247094 397024
rect 247052 396681 247080 397015
rect 247038 396672 247094 396681
rect 247038 396607 247094 396616
rect 246948 393984 247000 393990
rect 246948 393926 247000 393932
rect 246764 389904 246816 389910
rect 246764 389846 246816 389852
rect 246500 389146 246620 389174
rect 246592 352646 246620 389146
rect 246580 352640 246632 352646
rect 246580 352582 246632 352588
rect 246212 86284 246264 86290
rect 246212 86226 246264 86232
rect 246120 24472 246172 24478
rect 246120 24414 246172 24420
rect 246028 22772 246080 22778
rect 246028 22714 246080 22720
rect 246960 14754 246988 393926
rect 247144 392170 247172 400044
rect 247236 393786 247264 400044
rect 247328 398585 247356 400044
rect 247314 398576 247370 398585
rect 247314 398511 247370 398520
rect 247314 398304 247370 398313
rect 247314 398239 247370 398248
rect 247328 395622 247356 398239
rect 247316 395616 247368 395622
rect 247316 395558 247368 395564
rect 247224 393780 247276 393786
rect 247224 393722 247276 393728
rect 247420 393666 247448 400044
rect 247052 392142 247172 392170
rect 247236 393638 247448 393666
rect 246948 14748 247000 14754
rect 246948 14690 247000 14696
rect 245844 14680 245896 14686
rect 245844 14622 245896 14628
rect 247052 14618 247080 392142
rect 247132 392080 247184 392086
rect 247132 392022 247184 392028
rect 247040 14612 247092 14618
rect 247040 14554 247092 14560
rect 247144 14482 247172 392022
rect 247236 14550 247264 393638
rect 247316 393576 247368 393582
rect 247316 393518 247368 393524
rect 247328 24410 247356 393518
rect 247512 392170 247540 400044
rect 247604 398018 247632 400044
rect 247696 398138 247724 400044
rect 247684 398132 247736 398138
rect 247684 398074 247736 398080
rect 247604 397990 247724 398018
rect 247696 397254 247724 397990
rect 247592 397248 247644 397254
rect 247592 397190 247644 397196
rect 247684 397248 247736 397254
rect 247684 397190 247736 397196
rect 247420 392142 247540 392170
rect 247316 24404 247368 24410
rect 247316 24346 247368 24352
rect 247420 24342 247448 392142
rect 247500 392080 247552 392086
rect 247500 392022 247552 392028
rect 247408 24336 247460 24342
rect 247408 24278 247460 24284
rect 247512 24274 247540 392022
rect 247604 26926 247632 397190
rect 247684 395616 247736 395622
rect 247684 395558 247736 395564
rect 247696 393106 247724 395558
rect 247684 393100 247736 393106
rect 247684 393042 247736 393048
rect 247788 392154 247816 400044
rect 247776 392148 247828 392154
rect 247776 392090 247828 392096
rect 247880 392086 247908 400044
rect 247972 398313 248000 400044
rect 247958 398304 248014 398313
rect 247958 398239 248014 398248
rect 247960 398132 248012 398138
rect 247960 398074 248012 398080
rect 247972 394670 248000 398074
rect 248064 397497 248092 400044
rect 248156 397905 248184 400044
rect 248142 397896 248198 397905
rect 248142 397831 248198 397840
rect 248248 397769 248276 400044
rect 248234 397760 248290 397769
rect 248234 397695 248290 397704
rect 248340 397633 248368 400044
rect 248326 397624 248382 397633
rect 248326 397559 248382 397568
rect 248050 397488 248106 397497
rect 248050 397423 248106 397432
rect 247960 394664 248012 394670
rect 247960 394606 248012 394612
rect 248432 392086 248460 400044
rect 248524 398721 248552 400044
rect 248510 398712 248566 398721
rect 248510 398647 248566 398656
rect 248510 398440 248566 398449
rect 248510 398375 248566 398384
rect 248524 392698 248552 398375
rect 248512 392692 248564 392698
rect 248512 392634 248564 392640
rect 248616 392170 248644 400044
rect 248708 393650 248736 400044
rect 248800 398313 248828 400044
rect 248786 398304 248842 398313
rect 248786 398239 248842 398248
rect 248786 398168 248842 398177
rect 248786 398103 248842 398112
rect 248800 397594 248828 398103
rect 248788 397588 248840 397594
rect 248788 397530 248840 397536
rect 248696 393644 248748 393650
rect 248696 393586 248748 393592
rect 248892 392306 248920 400044
rect 248524 392142 248644 392170
rect 248708 392278 248920 392306
rect 247868 392080 247920 392086
rect 247868 392022 247920 392028
rect 248420 392080 248472 392086
rect 248420 392022 248472 392028
rect 248420 391944 248472 391950
rect 248420 391886 248472 391892
rect 247592 26920 247644 26926
rect 247592 26862 247644 26868
rect 247500 24268 247552 24274
rect 247500 24210 247552 24216
rect 247224 14544 247276 14550
rect 247224 14486 247276 14492
rect 247132 14476 247184 14482
rect 247132 14418 247184 14424
rect 245660 13116 245712 13122
rect 245660 13058 245712 13064
rect 243084 11824 243136 11830
rect 243084 11766 243136 11772
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 247592 4888 247644 4894
rect 247592 4830 247644 4836
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 242898 3496 242954 3505
rect 242898 3431 242954 3440
rect 242164 3188 242216 3194
rect 242164 3130 242216 3136
rect 242912 480 242940 3431
rect 244108 480 244136 3538
rect 246396 3392 246448 3398
rect 246396 3334 246448 3340
rect 245200 3188 245252 3194
rect 245200 3130 245252 3136
rect 245212 480 245240 3130
rect 246408 480 246436 3334
rect 247604 480 247632 4830
rect 248432 3602 248460 391886
rect 248524 7682 248552 392142
rect 248708 392034 248736 392278
rect 248788 392216 248840 392222
rect 248984 392170 249012 400044
rect 249076 398449 249104 400044
rect 249062 398440 249118 398449
rect 249062 398375 249118 398384
rect 249064 398336 249116 398342
rect 249064 398278 249116 398284
rect 249076 397730 249104 398278
rect 249064 397724 249116 397730
rect 249064 397666 249116 397672
rect 249064 397180 249116 397186
rect 249064 397122 249116 397128
rect 249076 396846 249104 397122
rect 249064 396840 249116 396846
rect 249064 396782 249116 396788
rect 248788 392158 248840 392164
rect 248616 392006 248736 392034
rect 248616 16250 248644 392006
rect 248696 391740 248748 391746
rect 248696 391682 248748 391688
rect 248604 16244 248656 16250
rect 248604 16186 248656 16192
rect 248708 16182 248736 391682
rect 248696 16176 248748 16182
rect 248696 16118 248748 16124
rect 248800 16114 248828 392158
rect 248892 392142 249012 392170
rect 248892 24138 248920 392142
rect 248972 392080 249024 392086
rect 248972 392022 249024 392028
rect 248984 24206 249012 392022
rect 249168 391746 249196 400044
rect 249156 391740 249208 391746
rect 249156 391682 249208 391688
rect 249260 389174 249288 400044
rect 249352 391950 249380 400044
rect 249444 392222 249472 400044
rect 249536 397633 249564 400044
rect 249522 397624 249578 397633
rect 249522 397559 249578 397568
rect 249628 397497 249656 400044
rect 249720 397769 249748 400044
rect 249706 397760 249762 397769
rect 249706 397695 249762 397704
rect 249614 397488 249670 397497
rect 249614 397423 249670 397432
rect 249432 392216 249484 392222
rect 249432 392158 249484 392164
rect 249340 391944 249392 391950
rect 249340 391886 249392 391892
rect 249812 389774 249840 400044
rect 249904 398177 249932 400044
rect 249890 398168 249946 398177
rect 249890 398103 249946 398112
rect 249996 392306 250024 400044
rect 250088 393938 250116 400044
rect 250180 395622 250208 400044
rect 250168 395616 250220 395622
rect 250168 395558 250220 395564
rect 250088 393910 250208 393938
rect 250076 393848 250128 393854
rect 250076 393790 250128 393796
rect 249904 392278 250024 392306
rect 249800 389768 249852 389774
rect 249800 389710 249852 389716
rect 249800 389632 249852 389638
rect 249800 389574 249852 389580
rect 249076 389146 249288 389174
rect 249076 82142 249104 389146
rect 249064 82136 249116 82142
rect 249064 82078 249116 82084
rect 249064 46232 249116 46238
rect 249064 46174 249116 46180
rect 248972 24200 249024 24206
rect 248972 24142 249024 24148
rect 248880 24132 248932 24138
rect 248880 24074 248932 24080
rect 248788 16108 248840 16114
rect 248788 16050 248840 16056
rect 248512 7676 248564 7682
rect 248512 7618 248564 7624
rect 249076 6914 249104 46174
rect 248800 6886 249104 6914
rect 248420 3596 248472 3602
rect 248420 3538 248472 3544
rect 248800 480 248828 6886
rect 249812 5166 249840 389574
rect 249904 16046 249932 392278
rect 249984 392216 250036 392222
rect 249984 392158 250036 392164
rect 249892 16040 249944 16046
rect 249892 15982 249944 15988
rect 249996 15910 250024 392158
rect 250088 15978 250116 393790
rect 250180 389858 250208 393910
rect 250272 393854 250300 400044
rect 250260 393848 250312 393854
rect 250260 393790 250312 393796
rect 250180 389830 250300 389858
rect 250168 389768 250220 389774
rect 250168 389710 250220 389716
rect 250180 355502 250208 389710
rect 250168 355496 250220 355502
rect 250168 355438 250220 355444
rect 250272 355434 250300 389830
rect 250364 356862 250392 400044
rect 250456 396030 250484 400044
rect 250444 396024 250496 396030
rect 250444 395966 250496 395972
rect 250444 395616 250496 395622
rect 250444 395558 250496 395564
rect 250456 392630 250484 395558
rect 250444 392624 250496 392630
rect 250444 392566 250496 392572
rect 250548 392222 250576 400044
rect 250536 392216 250588 392222
rect 250536 392158 250588 392164
rect 250444 391264 250496 391270
rect 250444 391206 250496 391212
rect 250352 356856 250404 356862
rect 250352 356798 250404 356804
rect 250260 355428 250312 355434
rect 250260 355370 250312 355376
rect 250076 15972 250128 15978
rect 250076 15914 250128 15920
rect 249984 15904 250036 15910
rect 249984 15846 250036 15852
rect 249800 5160 249852 5166
rect 249800 5102 249852 5108
rect 250456 3534 250484 391206
rect 250640 389174 250668 400044
rect 250732 389638 250760 400044
rect 250824 397633 250852 400044
rect 250810 397624 250866 397633
rect 250810 397559 250866 397568
rect 250916 396681 250944 400044
rect 251008 397497 251036 400044
rect 251100 397769 251128 400044
rect 251086 397760 251142 397769
rect 251086 397695 251142 397704
rect 250994 397488 251050 397497
rect 250994 397423 251050 397432
rect 250902 396672 250958 396681
rect 250902 396607 250958 396616
rect 250812 396024 250864 396030
rect 250812 395966 250864 395972
rect 250824 391338 250852 395966
rect 251192 393854 251220 400044
rect 251284 398041 251312 400044
rect 251270 398032 251326 398041
rect 251270 397967 251326 397976
rect 251272 394596 251324 394602
rect 251272 394538 251324 394544
rect 251180 393848 251232 393854
rect 251180 393790 251232 393796
rect 251180 393712 251232 393718
rect 251180 393654 251232 393660
rect 250812 391332 250864 391338
rect 250812 391274 250864 391280
rect 250720 389632 250772 389638
rect 250720 389574 250772 389580
rect 250548 389146 250668 389174
rect 250548 356794 250576 389146
rect 250536 356788 250588 356794
rect 250536 356730 250588 356736
rect 251192 4962 251220 393654
rect 251284 5030 251312 394538
rect 251376 393990 251404 400044
rect 251364 393984 251416 393990
rect 251364 393926 251416 393932
rect 251364 393848 251416 393854
rect 251364 393790 251416 393796
rect 251376 5098 251404 393790
rect 251468 7614 251496 400044
rect 251560 395078 251588 400044
rect 251548 395072 251600 395078
rect 251548 395014 251600 395020
rect 251548 393984 251600 393990
rect 251548 393926 251600 393932
rect 251652 393938 251680 400044
rect 251744 394074 251772 400044
rect 251836 394602 251864 400044
rect 251824 394596 251876 394602
rect 251824 394538 251876 394544
rect 251744 394046 251864 394074
rect 251560 17542 251588 393926
rect 251652 393910 251772 393938
rect 251640 393848 251692 393854
rect 251640 393790 251692 393796
rect 251548 17536 251600 17542
rect 251548 17478 251600 17484
rect 251652 17474 251680 393790
rect 251744 87650 251772 393910
rect 251836 356726 251864 394046
rect 251928 393854 251956 400044
rect 252020 395622 252048 400044
rect 252008 395616 252060 395622
rect 252008 395558 252060 395564
rect 252008 395072 252060 395078
rect 252008 395014 252060 395020
rect 251916 393848 251968 393854
rect 251916 393790 251968 393796
rect 252020 391270 252048 395014
rect 252112 393718 252140 400044
rect 252204 397769 252232 400044
rect 252190 397760 252246 397769
rect 252190 397695 252246 397704
rect 252296 397633 252324 400044
rect 252282 397624 252338 397633
rect 252282 397559 252338 397568
rect 252388 397497 252416 400044
rect 252480 397905 252508 400044
rect 252466 397896 252522 397905
rect 252466 397831 252522 397840
rect 252374 397488 252430 397497
rect 252374 397423 252430 397432
rect 252100 393712 252152 393718
rect 252100 393654 252152 393660
rect 252572 393038 252600 400044
rect 252664 398342 252692 400044
rect 252652 398336 252704 398342
rect 252652 398278 252704 398284
rect 252756 394058 252784 400044
rect 252744 394052 252796 394058
rect 252744 393994 252796 394000
rect 252848 393854 252876 400044
rect 252836 393848 252888 393854
rect 252836 393790 252888 393796
rect 252744 393780 252796 393786
rect 252744 393722 252796 393728
rect 252652 393712 252704 393718
rect 252652 393654 252704 393660
rect 252560 393032 252612 393038
rect 252560 392974 252612 392980
rect 252560 392760 252612 392766
rect 252560 392702 252612 392708
rect 252008 391264 252060 391270
rect 252008 391206 252060 391212
rect 251824 356720 251876 356726
rect 251824 356662 251876 356668
rect 251732 87644 251784 87650
rect 251732 87586 251784 87592
rect 251640 17468 251692 17474
rect 251640 17410 251692 17416
rect 251456 7608 251508 7614
rect 251456 7550 251508 7556
rect 251364 5092 251416 5098
rect 251364 5034 251416 5040
rect 251272 5024 251324 5030
rect 251272 4966 251324 4972
rect 251180 4956 251232 4962
rect 251180 4898 251232 4904
rect 252572 4826 252600 392702
rect 252664 4894 252692 393654
rect 252756 10334 252784 393722
rect 252940 393718 252968 400044
rect 252928 393712 252980 393718
rect 252928 393654 252980 393660
rect 253032 393394 253060 400044
rect 253124 395554 253152 400044
rect 253112 395548 253164 395554
rect 253112 395490 253164 395496
rect 253112 394052 253164 394058
rect 253112 393994 253164 394000
rect 252848 393366 253060 393394
rect 252848 17338 252876 393366
rect 252928 393304 252980 393310
rect 253124 393258 253152 393994
rect 253216 393938 253244 400044
rect 253308 394074 253336 400044
rect 253400 394176 253428 400044
rect 253492 394346 253520 400044
rect 253584 397633 253612 400044
rect 253676 399265 253704 400044
rect 253662 399256 253718 399265
rect 253662 399191 253718 399200
rect 253664 399084 253716 399090
rect 253664 399026 253716 399032
rect 253570 397624 253626 397633
rect 253570 397559 253626 397568
rect 253676 397526 253704 399026
rect 253664 397520 253716 397526
rect 253768 397497 253796 400044
rect 253860 397769 253888 400044
rect 253846 397760 253902 397769
rect 253846 397695 253902 397704
rect 253664 397462 253716 397468
rect 253754 397488 253810 397497
rect 253754 397423 253810 397432
rect 253952 395486 253980 400044
rect 254044 397526 254072 400044
rect 254032 397520 254084 397526
rect 254032 397462 254084 397468
rect 253940 395480 253992 395486
rect 253940 395422 253992 395428
rect 254136 394890 254164 400044
rect 254228 395418 254256 400044
rect 254320 398138 254348 400044
rect 254308 398132 254360 398138
rect 254308 398074 254360 398080
rect 254216 395412 254268 395418
rect 254216 395354 254268 395360
rect 254136 394862 254256 394890
rect 254032 394732 254084 394738
rect 254032 394674 254084 394680
rect 253940 394596 253992 394602
rect 253940 394538 253992 394544
rect 253492 394318 253612 394346
rect 253400 394148 253520 394176
rect 253308 394046 253428 394074
rect 253216 393910 253336 393938
rect 253204 393848 253256 393854
rect 253204 393790 253256 393796
rect 252928 393246 252980 393252
rect 252836 17332 252888 17338
rect 252836 17274 252888 17280
rect 252940 17270 252968 393246
rect 253032 393230 253152 393258
rect 253032 17406 253060 393230
rect 253216 393122 253244 393790
rect 253124 393094 253244 393122
rect 253124 354006 253152 393094
rect 253204 393032 253256 393038
rect 253204 392974 253256 392980
rect 253216 354074 253244 392974
rect 253308 355366 253336 393910
rect 253400 393310 253428 394046
rect 253492 393786 253520 394148
rect 253480 393780 253532 393786
rect 253480 393722 253532 393728
rect 253388 393304 253440 393310
rect 253388 393246 253440 393252
rect 253584 392766 253612 394318
rect 253664 393100 253716 393106
rect 253664 393042 253716 393048
rect 253676 392766 253704 393042
rect 253572 392760 253624 392766
rect 253572 392702 253624 392708
rect 253664 392760 253716 392766
rect 253664 392702 253716 392708
rect 253296 355360 253348 355366
rect 253296 355302 253348 355308
rect 253204 354068 253256 354074
rect 253204 354010 253256 354016
rect 253112 354000 253164 354006
rect 253112 353942 253164 353948
rect 253020 17400 253072 17406
rect 253020 17342 253072 17348
rect 252928 17264 252980 17270
rect 252928 17206 252980 17212
rect 252744 10328 252796 10334
rect 252744 10270 252796 10276
rect 253952 6254 253980 394538
rect 254044 6322 254072 394674
rect 254124 393916 254176 393922
rect 254124 393858 254176 393864
rect 254032 6316 254084 6322
rect 254032 6258 254084 6264
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254136 6186 254164 393858
rect 254228 18698 254256 394862
rect 254412 394738 254440 400044
rect 254400 394732 254452 394738
rect 254400 394674 254452 394680
rect 254504 394176 254532 400044
rect 254596 394602 254624 400044
rect 254584 394596 254636 394602
rect 254584 394538 254636 394544
rect 254412 394148 254532 394176
rect 254308 389428 254360 389434
rect 254308 389370 254360 389376
rect 254216 18692 254268 18698
rect 254216 18634 254268 18640
rect 254320 18630 254348 389370
rect 254412 25566 254440 394148
rect 254688 389434 254716 400044
rect 254780 395350 254808 400044
rect 254768 395344 254820 395350
rect 254768 395286 254820 395292
rect 254872 393922 254900 400044
rect 254860 393916 254912 393922
rect 254860 393858 254912 393864
rect 254676 389428 254728 389434
rect 254676 389370 254728 389376
rect 254964 389174 254992 400044
rect 255056 397633 255084 400044
rect 255042 397624 255098 397633
rect 255042 397559 255098 397568
rect 255148 397497 255176 400044
rect 255240 397769 255268 400044
rect 255226 397760 255282 397769
rect 255226 397695 255282 397704
rect 255134 397488 255190 397497
rect 255134 397423 255190 397432
rect 255226 395448 255282 395457
rect 255226 395383 255282 395392
rect 255240 394074 255268 395383
rect 255332 394176 255360 400044
rect 255424 398449 255452 400044
rect 255516 398682 255544 400044
rect 255504 398676 255556 398682
rect 255504 398618 255556 398624
rect 255410 398440 255466 398449
rect 255608 398410 255636 400044
rect 256056 399016 256108 399022
rect 256056 398958 256108 398964
rect 256068 398750 256096 398958
rect 263600 398880 263652 398886
rect 263600 398822 263652 398828
rect 256056 398744 256108 398750
rect 255962 398712 256018 398721
rect 256056 398686 256108 398692
rect 255962 398647 256018 398656
rect 255410 398375 255466 398384
rect 255596 398404 255648 398410
rect 255596 398346 255648 398352
rect 255332 394148 255452 394176
rect 255240 394046 255360 394074
rect 254504 389146 254992 389174
rect 254504 348430 254532 389146
rect 254492 348424 254544 348430
rect 254492 348366 254544 348372
rect 254400 25560 254452 25566
rect 254400 25502 254452 25508
rect 254308 18624 254360 18630
rect 254308 18566 254360 18572
rect 255332 16574 255360 394046
rect 255424 19990 255452 394148
rect 255412 19984 255464 19990
rect 255412 19926 255464 19932
rect 255332 16546 255912 16574
rect 254124 6180 254176 6186
rect 254124 6122 254176 6128
rect 254674 5264 254730 5273
rect 254674 5199 254730 5208
rect 252652 4888 252704 4894
rect 252652 4830 252704 4836
rect 252376 4820 252428 4826
rect 252376 4762 252428 4768
rect 252560 4820 252612 4826
rect 252560 4762 252612 4768
rect 250444 3528 250496 3534
rect 250444 3470 250496 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 249984 3392 250036 3398
rect 249984 3334 250036 3340
rect 249996 480 250024 3334
rect 251192 480 251220 3470
rect 252388 480 252416 4762
rect 253480 3460 253532 3466
rect 253480 3402 253532 3408
rect 253492 480 253520 3402
rect 254688 480 254716 5199
rect 255884 480 255912 16546
rect 255976 3534 256004 398647
rect 261484 398608 261536 398614
rect 261484 398550 261536 398556
rect 257528 398336 257580 398342
rect 257528 398278 257580 398284
rect 256700 398268 256752 398274
rect 256700 398210 256752 398216
rect 256424 397860 256476 397866
rect 256424 397802 256476 397808
rect 256332 397520 256384 397526
rect 256332 397462 256384 397468
rect 256148 397248 256200 397254
rect 256148 397190 256200 397196
rect 256056 397180 256108 397186
rect 256056 397122 256108 397128
rect 256068 3806 256096 397122
rect 256056 3800 256108 3806
rect 256056 3742 256108 3748
rect 256160 3602 256188 397190
rect 256240 395956 256292 395962
rect 256240 395898 256292 395904
rect 256252 4146 256280 395898
rect 256344 6390 256372 397462
rect 256436 27062 256464 397802
rect 256608 397792 256660 397798
rect 256608 397734 256660 397740
rect 256516 397724 256568 397730
rect 256516 397666 256568 397672
rect 256528 27130 256556 397666
rect 256620 83570 256648 397734
rect 256608 83564 256660 83570
rect 256608 83506 256660 83512
rect 256516 27124 256568 27130
rect 256516 27066 256568 27072
rect 256424 27056 256476 27062
rect 256424 26998 256476 27004
rect 256332 6384 256384 6390
rect 256332 6326 256384 6332
rect 256240 4140 256292 4146
rect 256240 4082 256292 4088
rect 256148 3596 256200 3602
rect 256148 3538 256200 3544
rect 255964 3528 256016 3534
rect 255964 3470 256016 3476
rect 256712 3398 256740 398210
rect 257436 397588 257488 397594
rect 257436 397530 257488 397536
rect 257342 395584 257398 395593
rect 257342 395519 257398 395528
rect 257356 3738 257384 395519
rect 257448 12102 257476 397530
rect 257540 71738 257568 398278
rect 259552 398064 259604 398070
rect 259552 398006 259604 398012
rect 258816 397996 258868 398002
rect 258816 397938 258868 397944
rect 257620 397656 257672 397662
rect 257620 397598 257672 397604
rect 257632 334626 257660 397598
rect 258724 394664 258776 394670
rect 258724 394606 258776 394612
rect 257620 334620 257672 334626
rect 257620 334562 257672 334568
rect 257528 71732 257580 71738
rect 257528 71674 257580 71680
rect 257436 12096 257488 12102
rect 257436 12038 257488 12044
rect 257344 3732 257396 3738
rect 257344 3674 257396 3680
rect 258736 3670 258764 394606
rect 258828 305658 258856 397938
rect 258816 305652 258868 305658
rect 258816 305594 258868 305600
rect 259564 16574 259592 398006
rect 260102 397896 260158 397905
rect 260102 397831 260158 397840
rect 260116 336054 260144 397831
rect 260104 336048 260156 336054
rect 260104 335990 260156 335996
rect 261496 186998 261524 398550
rect 261484 186992 261536 186998
rect 261484 186934 261536 186940
rect 263612 16574 263640 398822
rect 264244 398540 264296 398546
rect 264244 398482 264296 398488
rect 264256 29646 264284 398482
rect 264336 398472 264388 398478
rect 264336 398414 264388 398420
rect 264348 188358 264376 398414
rect 264992 398342 265020 446655
rect 282380 446282 282408 580246
rect 282932 463214 282960 702406
rect 300136 700534 300164 703520
rect 296076 700528 296128 700534
rect 296076 700470 296128 700476
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 293224 700460 293276 700466
rect 293224 700402 293276 700408
rect 291844 700392 291896 700398
rect 291844 700334 291896 700340
rect 286324 696992 286376 696998
rect 286324 696934 286376 696940
rect 284300 597304 284352 597310
rect 284300 597246 284352 597252
rect 284312 596698 284340 597246
rect 284576 596896 284628 596902
rect 284576 596838 284628 596844
rect 284392 596828 284444 596834
rect 284392 596770 284444 596776
rect 284300 596692 284352 596698
rect 284300 596634 284352 596640
rect 283104 596624 283156 596630
rect 283104 596566 283156 596572
rect 283012 596556 283064 596562
rect 283012 596498 283064 596504
rect 282920 463208 282972 463214
rect 282920 463150 282972 463156
rect 283024 452334 283052 596498
rect 283116 596358 283144 596566
rect 283104 596352 283156 596358
rect 283104 596294 283156 596300
rect 283012 452328 283064 452334
rect 283012 452270 283064 452276
rect 283116 452130 283144 596294
rect 283564 583024 283616 583030
rect 283564 582966 283616 582972
rect 283104 452124 283156 452130
rect 283104 452066 283156 452072
rect 283576 447030 283604 582966
rect 284312 452538 284340 596634
rect 284404 596290 284432 596770
rect 284588 596494 284616 596838
rect 284484 596488 284536 596494
rect 284484 596430 284536 596436
rect 284576 596488 284628 596494
rect 284576 596430 284628 596436
rect 284496 596358 284524 596430
rect 284484 596352 284536 596358
rect 284484 596294 284536 596300
rect 284392 596284 284444 596290
rect 284392 596226 284444 596232
rect 284300 452532 284352 452538
rect 284300 452474 284352 452480
rect 284404 452470 284432 596226
rect 284392 452464 284444 452470
rect 284392 452406 284444 452412
rect 284496 452402 284524 596294
rect 284484 452396 284536 452402
rect 284484 452338 284536 452344
rect 284588 452266 284616 596430
rect 284944 590708 284996 590714
rect 284944 590650 284996 590656
rect 284956 453422 284984 590650
rect 285036 580372 285088 580378
rect 285036 580314 285088 580320
rect 284944 453416 284996 453422
rect 284944 453358 284996 453364
rect 284576 452260 284628 452266
rect 284576 452202 284628 452208
rect 283564 447024 283616 447030
rect 283564 446966 283616 446972
rect 285048 446894 285076 580314
rect 286336 451926 286364 696934
rect 289084 589960 289136 589966
rect 289084 589902 289136 589908
rect 287704 588668 287756 588674
rect 287704 588610 287756 588616
rect 286416 587172 286468 587178
rect 286416 587114 286468 587120
rect 286324 451920 286376 451926
rect 286324 451862 286376 451868
rect 285036 446888 285088 446894
rect 285036 446830 285088 446836
rect 286428 446350 286456 587114
rect 287716 446690 287744 588610
rect 287796 498840 287848 498846
rect 287796 498782 287848 498788
rect 287808 488034 287836 498782
rect 287796 488028 287848 488034
rect 287796 487970 287848 487976
rect 287704 446684 287756 446690
rect 287704 446626 287756 446632
rect 289096 446622 289124 589902
rect 289176 581664 289228 581670
rect 289176 581606 289228 581612
rect 289188 446826 289216 581606
rect 291856 461854 291884 700334
rect 291936 488436 291988 488442
rect 291936 488378 291988 488384
rect 291844 461848 291896 461854
rect 291844 461790 291896 461796
rect 291948 449585 291976 488378
rect 293236 460358 293264 700402
rect 295984 700324 296036 700330
rect 295984 700266 296036 700272
rect 293316 584452 293368 584458
rect 293316 584394 293368 584400
rect 293224 460352 293276 460358
rect 293224 460294 293276 460300
rect 293224 458312 293276 458318
rect 293224 458254 293276 458260
rect 293236 450838 293264 458254
rect 293224 450832 293276 450838
rect 293224 450774 293276 450780
rect 291934 449576 291990 449585
rect 291934 449511 291990 449520
rect 293224 448860 293276 448866
rect 293224 448802 293276 448808
rect 293132 447364 293184 447370
rect 293132 447306 293184 447312
rect 289176 446820 289228 446826
rect 289176 446762 289228 446768
rect 289084 446616 289136 446622
rect 289084 446558 289136 446564
rect 286416 446344 286468 446350
rect 286416 446286 286468 446292
rect 282368 446276 282420 446282
rect 282368 446218 282420 446224
rect 266176 445528 266228 445534
rect 266176 445470 266228 445476
rect 265806 444952 265862 444961
rect 265806 444887 265862 444896
rect 265622 444816 265678 444825
rect 265622 444751 265678 444760
rect 265532 443148 265584 443154
rect 265532 443090 265584 443096
rect 265544 436082 265572 443090
rect 265532 436076 265584 436082
rect 265532 436018 265584 436024
rect 264980 398336 265032 398342
rect 264980 398278 265032 398284
rect 264992 397934 265020 398278
rect 264980 397928 265032 397934
rect 264980 397870 265032 397876
rect 264336 188352 264388 188358
rect 264336 188294 264388 188300
rect 265636 46918 265664 444751
rect 265714 443456 265770 443465
rect 265714 443391 265770 443400
rect 265728 73166 265756 443391
rect 265820 86970 265848 444887
rect 266084 444440 266136 444446
rect 266084 444382 266136 444388
rect 265898 443728 265954 443737
rect 265898 443663 265954 443672
rect 265912 139398 265940 443663
rect 265992 443420 266044 443426
rect 265992 443362 266044 443368
rect 266004 299470 266032 443362
rect 266096 398002 266124 444382
rect 266188 404326 266216 445470
rect 273904 445324 273956 445330
rect 273904 445266 273956 445272
rect 269856 445188 269908 445194
rect 269856 445130 269908 445136
rect 268476 445120 268528 445126
rect 268476 445062 268528 445068
rect 267096 444984 267148 444990
rect 267096 444926 267148 444932
rect 266360 443284 266412 443290
rect 266360 443226 266412 443232
rect 266372 440230 266400 443226
rect 267004 443080 267056 443086
rect 267004 443022 267056 443028
rect 266360 440224 266412 440230
rect 266360 440166 266412 440172
rect 267016 408474 267044 443022
rect 267108 431934 267136 444926
rect 268384 444848 268436 444854
rect 268384 444790 268436 444796
rect 267096 431928 267148 431934
rect 267096 431870 267148 431876
rect 267004 408468 267056 408474
rect 267004 408410 267056 408416
rect 266176 404320 266228 404326
rect 266176 404262 266228 404268
rect 266084 397996 266136 398002
rect 266084 397938 266136 397944
rect 266360 395888 266412 395894
rect 266360 395830 266412 395836
rect 265992 299464 266044 299470
rect 265992 299406 266044 299412
rect 265900 139392 265952 139398
rect 265900 139334 265952 139340
rect 265808 86964 265860 86970
rect 265808 86906 265860 86912
rect 265716 73160 265768 73166
rect 265716 73102 265768 73108
rect 265624 46912 265676 46918
rect 265624 46854 265676 46860
rect 264244 29640 264296 29646
rect 264244 29582 264296 29588
rect 266372 16574 266400 395830
rect 267740 392964 267792 392970
rect 267740 392906 267792 392912
rect 259564 16546 260696 16574
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 259460 4140 259512 4146
rect 259460 4082 259512 4088
rect 258264 3664 258316 3670
rect 258264 3606 258316 3612
rect 258724 3664 258776 3670
rect 258724 3606 258776 3612
rect 256700 3392 256752 3398
rect 256700 3334 256752 3340
rect 257066 3360 257122 3369
rect 257066 3295 257122 3304
rect 257080 480 257108 3295
rect 258276 480 258304 3606
rect 259472 480 259500 4082
rect 260668 480 260696 16546
rect 262956 5228 263008 5234
rect 262956 5170 263008 5176
rect 261760 3868 261812 3874
rect 261760 3810 261812 3816
rect 261772 480 261800 3810
rect 262968 480 262996 5170
rect 264164 480 264192 16546
rect 264980 12232 265032 12238
rect 264980 12174 265032 12180
rect 221526 354 221638 480
rect 221384 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 12174
rect 266556 480 266584 16546
rect 267752 480 267780 392906
rect 268396 245614 268424 444790
rect 268488 426426 268516 445062
rect 268476 426420 268528 426426
rect 268476 426362 268528 426368
rect 269764 398676 269816 398682
rect 269764 398618 269816 398624
rect 269120 395820 269172 395826
rect 269120 395762 269172 395768
rect 268384 245608 268436 245614
rect 268384 245550 268436 245556
rect 267832 19168 267884 19174
rect 267832 19110 267884 19116
rect 267844 16574 267872 19110
rect 269132 16574 269160 395762
rect 269776 167686 269804 398618
rect 269868 353258 269896 445130
rect 271142 398576 271198 398585
rect 271142 398511 271198 398520
rect 269856 353252 269908 353258
rect 269856 353194 269908 353200
rect 270500 352912 270552 352918
rect 270500 352854 270552 352860
rect 269764 167680 269816 167686
rect 269764 167622 269816 167628
rect 270512 16574 270540 352854
rect 271156 31074 271184 398511
rect 273258 177304 273314 177313
rect 273258 177239 273314 177248
rect 271144 31068 271196 31074
rect 271144 31010 271196 31016
rect 271880 19100 271932 19106
rect 271880 19042 271932 19048
rect 271892 16574 271920 19042
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 177239
rect 273916 126954 273944 445266
rect 275284 444780 275336 444786
rect 275284 444722 275336 444728
rect 275296 167006 275324 444722
rect 278044 444712 278096 444718
rect 278044 444654 278096 444660
rect 283562 444680 283618 444689
rect 277400 399084 277452 399090
rect 277400 399026 277452 399032
rect 275376 398404 275428 398410
rect 275376 398346 275428 398352
rect 275388 191146 275416 398346
rect 276020 395752 276072 395758
rect 276020 395694 276072 395700
rect 275376 191140 275428 191146
rect 275376 191082 275428 191088
rect 275284 167000 275336 167006
rect 275284 166942 275336 166948
rect 273904 126948 273956 126954
rect 273904 126890 273956 126896
rect 274822 6488 274878 6497
rect 274822 6423 274878 6432
rect 274836 480 274864 6423
rect 276032 3874 276060 395694
rect 276110 18592 276166 18601
rect 276110 18527 276166 18536
rect 276020 3868 276072 3874
rect 276020 3810 276072 3816
rect 276124 3482 276152 18527
rect 277412 16574 277440 399026
rect 278056 153202 278084 444654
rect 283562 444615 283618 444624
rect 281540 355632 281592 355638
rect 281540 355574 281592 355580
rect 278044 153196 278096 153202
rect 278044 153138 278096 153144
rect 280160 25968 280212 25974
rect 280160 25910 280212 25916
rect 278780 19032 278832 19038
rect 278780 18974 278832 18980
rect 278792 16574 278820 18974
rect 280172 16574 280200 25910
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276756 3868 276808 3874
rect 276756 3810 276808 3816
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3810
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 355574
rect 283576 60722 283604 444615
rect 292946 442776 293002 442785
rect 292946 442711 293002 442720
rect 292960 400897 292988 442711
rect 293144 401033 293172 447306
rect 293130 401024 293186 401033
rect 293130 400959 293186 400968
rect 292946 400888 293002 400897
rect 292946 400823 293002 400832
rect 293236 398614 293264 448802
rect 293328 446758 293356 584394
rect 293868 527060 293920 527066
rect 293868 527002 293920 527008
rect 293880 489914 293908 527002
rect 293420 489886 293908 489914
rect 293420 488073 293448 489886
rect 293406 488064 293462 488073
rect 293406 487999 293462 488008
rect 293420 477494 293448 487999
rect 293408 477488 293460 477494
rect 293408 477430 293460 477436
rect 295996 454714 296024 700266
rect 296088 468654 296116 700470
rect 332520 700466 332548 703520
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364996 700330 365024 703520
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 397472 699718 397500 703520
rect 413664 700602 413692 703520
rect 405004 700596 405056 700602
rect 405004 700538 405056 700544
rect 413652 700596 413704 700602
rect 413652 700538 413704 700544
rect 403624 700460 403676 700466
rect 403624 700402 403676 700408
rect 399484 700392 399536 700398
rect 399484 700334 399536 700340
rect 395344 699712 395396 699718
rect 395344 699654 395396 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 297914 636984 297970 636993
rect 297914 636919 297970 636928
rect 297822 634264 297878 634273
rect 297822 634199 297878 634208
rect 297638 633176 297694 633185
rect 297638 633111 297694 633120
rect 297454 631544 297510 631553
rect 297454 631479 297510 631488
rect 296994 610192 297050 610201
rect 296994 610127 297050 610136
rect 296902 608288 296958 608297
rect 296902 608223 296958 608232
rect 296810 521520 296866 521529
rect 296810 521455 296866 521464
rect 296824 488345 296852 521455
rect 296916 498273 296944 608223
rect 297008 500857 297036 610127
rect 297086 608696 297142 608705
rect 297086 608631 297142 608640
rect 296994 500848 297050 500857
rect 296994 500783 297050 500792
rect 297100 498846 297128 608631
rect 297364 600296 297416 600302
rect 297364 600238 297416 600244
rect 297272 598052 297324 598058
rect 297272 597994 297324 598000
rect 297180 585200 297232 585206
rect 297180 585142 297232 585148
rect 297192 526017 297220 585142
rect 297284 527066 297312 597994
rect 297272 527060 297324 527066
rect 297272 527002 297324 527008
rect 297178 526008 297234 526017
rect 297178 525943 297234 525952
rect 297088 498840 297140 498846
rect 297088 498782 297140 498788
rect 297100 498681 297128 498782
rect 297086 498672 297142 498681
rect 297086 498607 297142 498616
rect 296902 498264 296958 498273
rect 296902 498199 296958 498208
rect 296810 488336 296866 488345
rect 296810 488271 296866 488280
rect 296824 485994 296852 488271
rect 296812 485988 296864 485994
rect 296812 485930 296864 485936
rect 296076 468648 296128 468654
rect 296076 468590 296128 468596
rect 296076 458652 296128 458658
rect 296076 458594 296128 458600
rect 295984 454708 296036 454714
rect 295984 454650 296036 454656
rect 293592 448996 293644 449002
rect 293592 448938 293644 448944
rect 293408 448656 293460 448662
rect 293408 448598 293460 448604
rect 293316 446752 293368 446758
rect 293316 446694 293368 446700
rect 293316 444508 293368 444514
rect 293316 444450 293368 444456
rect 293328 400110 293356 444450
rect 293316 400104 293368 400110
rect 293316 400046 293368 400052
rect 293224 398608 293276 398614
rect 293224 398550 293276 398556
rect 293420 398070 293448 448598
rect 293500 447432 293552 447438
rect 293500 447374 293552 447380
rect 293512 398342 293540 447374
rect 293604 400994 293632 448938
rect 293684 448928 293736 448934
rect 293684 448870 293736 448876
rect 293592 400988 293644 400994
rect 293592 400930 293644 400936
rect 293696 400926 293724 448870
rect 293868 448792 293920 448798
rect 293868 448734 293920 448740
rect 293776 448588 293828 448594
rect 293776 448530 293828 448536
rect 293788 401062 293816 448530
rect 293880 401130 293908 448734
rect 296088 447846 296116 458594
rect 297192 449721 297220 525943
rect 297376 524385 297404 600238
rect 297468 598874 297496 631479
rect 297546 628552 297602 628561
rect 297546 628487 297602 628496
rect 297456 598868 297508 598874
rect 297456 598810 297508 598816
rect 297362 524376 297418 524385
rect 297362 524311 297418 524320
rect 297270 521656 297326 521665
rect 297270 521591 297326 521600
rect 297284 520305 297312 521591
rect 297270 520296 297326 520305
rect 297270 520231 297326 520240
rect 297284 488374 297312 520231
rect 297376 489841 297404 524311
rect 297468 521529 297496 598810
rect 297560 598806 297588 628487
rect 297548 598800 297600 598806
rect 297548 598742 297600 598748
rect 297454 521520 297510 521529
rect 297454 521455 297510 521464
rect 297560 518673 297588 598742
rect 297652 523297 297680 633111
rect 297730 630184 297786 630193
rect 297730 630119 297786 630128
rect 297638 523288 297694 523297
rect 297638 523223 297694 523232
rect 297546 518664 297602 518673
rect 297546 518599 297602 518608
rect 297560 517585 297588 518599
rect 297546 517576 297602 517585
rect 297546 517511 297602 517520
rect 297362 489832 297418 489841
rect 297652 489802 297680 523223
rect 297744 521665 297772 630119
rect 297836 600302 297864 634199
rect 297824 600296 297876 600302
rect 297824 600238 297876 600244
rect 297836 600030 297864 600238
rect 297824 600024 297876 600030
rect 297824 599966 297876 599972
rect 297928 598942 297956 636919
rect 298006 635896 298062 635905
rect 298006 635831 298062 635840
rect 297916 598936 297968 598942
rect 297916 598878 297968 598884
rect 297928 598058 297956 598878
rect 297916 598052 297968 598058
rect 297916 597994 297968 598000
rect 298020 585818 298048 635831
rect 318338 597544 318394 597553
rect 318338 597479 318394 597488
rect 319442 597544 319498 597553
rect 319442 597479 319498 597488
rect 320086 597544 320142 597553
rect 320086 597479 320142 597488
rect 320914 597544 320970 597553
rect 320914 597479 320970 597488
rect 322294 597544 322350 597553
rect 322294 597479 322350 597488
rect 322938 597544 322994 597553
rect 322938 597479 322994 597488
rect 324318 597544 324374 597553
rect 324318 597479 324374 597488
rect 325790 597544 325846 597553
rect 325790 597479 325846 597488
rect 329838 597544 329894 597553
rect 329838 597479 329894 597488
rect 345018 597544 345074 597553
rect 345018 597479 345074 597488
rect 360198 597544 360254 597553
rect 360198 597479 360254 597488
rect 318352 597174 318380 597479
rect 319456 597242 319484 597479
rect 319444 597236 319496 597242
rect 319444 597178 319496 597184
rect 318340 597168 318392 597174
rect 318340 597110 318392 597116
rect 314658 597000 314714 597009
rect 314658 596935 314714 596944
rect 313278 596864 313334 596873
rect 299204 596828 299256 596834
rect 313278 596799 313280 596808
rect 299204 596770 299256 596776
rect 313332 596799 313334 596808
rect 313280 596770 313332 596776
rect 298836 585880 298888 585886
rect 298836 585822 298888 585828
rect 298008 585812 298060 585818
rect 298008 585754 298060 585760
rect 298020 585206 298048 585754
rect 298008 585200 298060 585206
rect 298008 585142 298060 585148
rect 298006 527096 298062 527105
rect 298006 527031 298008 527040
rect 298060 527031 298062 527040
rect 298008 527002 298060 527008
rect 297730 521656 297786 521665
rect 297730 521591 297786 521600
rect 298006 517576 298062 517585
rect 298006 517511 298062 517520
rect 297914 500848 297970 500857
rect 297914 500783 297970 500792
rect 297928 500313 297956 500783
rect 297914 500304 297970 500313
rect 297914 500239 297970 500248
rect 297822 498264 297878 498273
rect 297822 498199 297878 498208
rect 297362 489767 297418 489776
rect 297640 489796 297692 489802
rect 297272 488368 297324 488374
rect 297272 488310 297324 488316
rect 297284 486062 297312 488310
rect 297272 486056 297324 486062
rect 297272 485998 297324 486004
rect 297376 449857 297404 489767
rect 297640 489738 297692 489744
rect 297652 486690 297680 489738
rect 297836 488442 297864 498199
rect 297824 488436 297876 488442
rect 297824 488378 297876 488384
rect 297928 488170 297956 500239
rect 298020 488209 298048 517511
rect 298006 488200 298062 488209
rect 297916 488164 297968 488170
rect 298006 488135 298062 488144
rect 297916 488106 297968 488112
rect 297468 486662 297680 486690
rect 297362 449848 297418 449857
rect 297362 449783 297418 449792
rect 297178 449712 297234 449721
rect 297178 449647 297234 449656
rect 296536 448724 296588 448730
rect 296536 448666 296588 448672
rect 296076 447840 296128 447846
rect 296076 447782 296128 447788
rect 296260 447160 296312 447166
rect 296260 447102 296312 447108
rect 295892 445800 295944 445806
rect 295892 445742 295944 445748
rect 295800 443896 295852 443902
rect 295800 443838 295852 443844
rect 293868 401124 293920 401130
rect 293868 401066 293920 401072
rect 293776 401056 293828 401062
rect 293776 400998 293828 401004
rect 293684 400920 293736 400926
rect 293684 400862 293736 400868
rect 295812 398410 295840 443838
rect 295904 398750 295932 445742
rect 296074 444544 296130 444553
rect 296074 444479 296130 444488
rect 295982 442368 296038 442377
rect 295982 442303 296038 442312
rect 295892 398744 295944 398750
rect 295892 398686 295944 398692
rect 295800 398404 295852 398410
rect 295800 398346 295852 398352
rect 293500 398336 293552 398342
rect 293500 398278 293552 398284
rect 293408 398064 293460 398070
rect 293408 398006 293460 398012
rect 291198 393952 291254 393961
rect 291198 393887 291254 393896
rect 288440 355564 288492 355570
rect 288440 355506 288492 355512
rect 287060 87780 287112 87786
rect 287060 87722 287112 87728
rect 283564 60716 283616 60722
rect 283564 60658 283616 60664
rect 284300 25900 284352 25906
rect 284300 25842 284352 25848
rect 282920 18964 282972 18970
rect 282920 18906 282972 18912
rect 282932 16574 282960 18906
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 25842
rect 285680 20256 285732 20262
rect 285680 20198 285732 20204
rect 285692 16574 285720 20198
rect 287072 16574 287100 87722
rect 288452 16574 288480 355506
rect 289818 20224 289874 20233
rect 289818 20159 289874 20168
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 285404 6520 285456 6526
rect 285404 6462 285456 6468
rect 285416 480 285444 6462
rect 286612 480 286640 16546
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 20159
rect 291212 16574 291240 393887
rect 295340 392896 295392 392902
rect 295340 392838 295392 392844
rect 293960 390040 294012 390046
rect 293960 389982 294012 389988
rect 292578 20088 292634 20097
rect 292578 20023 292634 20032
rect 292592 16574 292620 20023
rect 293972 16574 294000 389982
rect 295352 16574 295380 392838
rect 295996 179382 296024 442303
rect 295984 179376 296036 179382
rect 295984 179318 296036 179324
rect 296088 100706 296116 444479
rect 296166 442232 296222 442241
rect 296166 442167 296222 442176
rect 296180 219434 296208 442167
rect 296272 313274 296300 447102
rect 296444 444644 296496 444650
rect 296444 444586 296496 444592
rect 296350 442504 296406 442513
rect 296350 442439 296406 442448
rect 296260 313268 296312 313274
rect 296260 313210 296312 313216
rect 296364 259418 296392 442439
rect 296456 365702 296484 444586
rect 296548 398478 296576 448666
rect 297468 448322 297496 486662
rect 297928 486282 297956 488106
rect 297560 486254 297956 486282
rect 297456 448316 297508 448322
rect 297456 448258 297508 448264
rect 297560 448254 297588 486254
rect 298020 486146 298048 488135
rect 297652 486118 298048 486146
rect 297652 448526 297680 486118
rect 297732 486056 297784 486062
rect 297732 485998 297784 486004
rect 297640 448520 297692 448526
rect 297640 448462 297692 448468
rect 297744 448458 297772 485998
rect 297916 485988 297968 485994
rect 297916 485930 297968 485936
rect 297822 452432 297878 452441
rect 297822 452367 297878 452376
rect 297836 451314 297864 452367
rect 297824 451308 297876 451314
rect 297824 451250 297876 451256
rect 297732 448452 297784 448458
rect 297732 448394 297784 448400
rect 297928 448390 297956 485930
rect 298744 458516 298796 458522
rect 298744 458458 298796 458464
rect 298008 458448 298060 458454
rect 298008 458390 298060 458396
rect 298020 450770 298048 458390
rect 298008 450764 298060 450770
rect 298008 450706 298060 450712
rect 298756 449274 298784 458458
rect 298744 449268 298796 449274
rect 298744 449210 298796 449216
rect 297916 448384 297968 448390
rect 297916 448326 297968 448332
rect 298006 448352 298062 448361
rect 298006 448287 298062 448296
rect 297548 448248 297600 448254
rect 297548 448190 297600 448196
rect 298020 447506 298048 448287
rect 298008 447500 298060 447506
rect 298008 447442 298060 447448
rect 296628 447296 296680 447302
rect 296628 447238 296680 447244
rect 296640 398818 296668 447238
rect 298652 447228 298704 447234
rect 298652 447170 298704 447176
rect 298100 446548 298152 446554
rect 298100 446490 298152 446496
rect 298112 446457 298140 446490
rect 298098 446448 298154 446457
rect 298098 446383 298154 446392
rect 297364 443828 297416 443834
rect 297364 443770 297416 443776
rect 297180 436076 297232 436082
rect 297180 436018 297232 436024
rect 297192 434761 297220 436018
rect 297178 434752 297234 434761
rect 297178 434687 297234 434696
rect 297376 413001 297404 443770
rect 297456 443760 297508 443766
rect 297456 443702 297508 443708
rect 297468 417081 297496 443702
rect 297548 443692 297600 443698
rect 297548 443634 297600 443640
rect 297560 421841 297588 443634
rect 298006 443592 298062 443601
rect 298006 443527 298062 443536
rect 298020 443018 298048 443527
rect 298560 443352 298612 443358
rect 298560 443294 298612 443300
rect 298008 443012 298060 443018
rect 298008 442954 298060 442960
rect 298008 440224 298060 440230
rect 298008 440166 298060 440172
rect 298020 439521 298048 440166
rect 298006 439512 298062 439521
rect 298006 439447 298062 439456
rect 298008 431928 298060 431934
rect 298008 431870 298060 431876
rect 298020 430681 298048 431870
rect 298006 430672 298062 430681
rect 298006 430607 298062 430616
rect 298008 426420 298060 426426
rect 298008 426362 298060 426368
rect 298020 425921 298048 426362
rect 298006 425912 298062 425921
rect 298006 425847 298062 425856
rect 297546 421832 297602 421841
rect 297546 421767 297602 421776
rect 297454 417072 297510 417081
rect 297454 417007 297510 417016
rect 297362 412992 297418 413001
rect 297362 412927 297418 412936
rect 298008 408468 298060 408474
rect 298008 408410 298060 408416
rect 298020 408241 298048 408410
rect 298006 408232 298062 408241
rect 298006 408167 298062 408176
rect 298008 404320 298060 404326
rect 298008 404262 298060 404268
rect 298020 404161 298048 404262
rect 298006 404152 298062 404161
rect 298006 404087 298062 404096
rect 298572 400178 298600 443294
rect 298560 400172 298612 400178
rect 298560 400114 298612 400120
rect 296628 398812 296680 398818
rect 296628 398754 296680 398760
rect 296536 398472 296588 398478
rect 296536 398414 296588 398420
rect 298664 398274 298692 447170
rect 298848 446418 298876 585822
rect 299216 488306 299244 596770
rect 314672 596698 314700 596935
rect 318352 596766 318380 597110
rect 319260 597100 319312 597106
rect 319260 597042 319312 597048
rect 318340 596760 318392 596766
rect 318340 596702 318392 596708
rect 299296 596692 299348 596698
rect 299296 596634 299348 596640
rect 314660 596692 314712 596698
rect 314660 596634 314712 596640
rect 299204 488300 299256 488306
rect 299204 488242 299256 488248
rect 299216 487898 299244 488242
rect 299308 488238 299336 596634
rect 319272 596630 319300 597042
rect 319260 596624 319312 596630
rect 311898 596592 311954 596601
rect 319260 596566 319312 596572
rect 311898 596527 311954 596536
rect 311912 596222 311940 596527
rect 319456 596426 319484 597178
rect 320100 597106 320128 597479
rect 320088 597100 320140 597106
rect 320088 597042 320140 597048
rect 320928 597038 320956 597479
rect 320916 597032 320968 597038
rect 320916 596974 320968 596980
rect 320928 596562 320956 596974
rect 322308 596902 322336 597479
rect 321560 596896 321612 596902
rect 321560 596838 321612 596844
rect 322296 596896 322348 596902
rect 322296 596838 322348 596844
rect 320916 596556 320968 596562
rect 320916 596498 320968 596504
rect 321572 596494 321600 596838
rect 322952 596834 322980 597479
rect 322940 596828 322992 596834
rect 322940 596770 322992 596776
rect 321560 596488 321612 596494
rect 321560 596430 321612 596436
rect 319444 596420 319496 596426
rect 319444 596362 319496 596368
rect 322952 596358 322980 596770
rect 322940 596352 322992 596358
rect 322940 596294 322992 596300
rect 299388 596216 299440 596222
rect 299388 596158 299440 596164
rect 311900 596216 311952 596222
rect 311900 596158 311952 596164
rect 299296 488232 299348 488238
rect 299296 488174 299348 488180
rect 299204 487892 299256 487898
rect 299204 487834 299256 487840
rect 299308 487830 299336 488174
rect 299296 487824 299348 487830
rect 299296 487766 299348 487772
rect 299400 487150 299428 596158
rect 324332 588674 324360 597479
rect 324410 597408 324466 597417
rect 324410 597343 324466 597352
rect 324424 596970 324452 597343
rect 325804 597310 325832 597479
rect 325792 597304 325844 597310
rect 325792 597246 325844 597252
rect 324412 596964 324464 596970
rect 324412 596906 324464 596912
rect 324424 596290 324452 596906
rect 324412 596284 324464 596290
rect 324412 596226 324464 596232
rect 329852 589966 329880 597479
rect 339498 597000 339554 597009
rect 339498 596935 339554 596944
rect 335358 596320 335414 596329
rect 335358 596255 335414 596264
rect 329840 589960 329892 589966
rect 329840 589902 329892 589908
rect 324320 588668 324372 588674
rect 324320 588610 324372 588616
rect 335372 580378 335400 596255
rect 339512 583030 339540 596935
rect 339500 583024 339552 583030
rect 339500 582966 339552 582972
rect 345032 581670 345060 597479
rect 349158 597136 349214 597145
rect 349158 597071 349214 597080
rect 349172 584458 349200 597071
rect 354678 596320 354734 596329
rect 354678 596255 354734 596264
rect 354692 585886 354720 596255
rect 360212 587178 360240 597479
rect 360200 587172 360252 587178
rect 360200 587114 360252 587120
rect 354680 585880 354732 585886
rect 354680 585822 354732 585828
rect 349160 584452 349212 584458
rect 349160 584394 349212 584400
rect 345020 581664 345072 581670
rect 345020 581606 345072 581612
rect 335360 580372 335412 580378
rect 335360 580314 335412 580320
rect 314290 488472 314346 488481
rect 314290 488407 314346 488416
rect 315394 488472 315450 488481
rect 315394 488407 315450 488416
rect 322938 488472 322994 488481
rect 322938 488407 322994 488416
rect 314304 488306 314332 488407
rect 314292 488300 314344 488306
rect 314292 488242 314344 488248
rect 315408 488238 315436 488407
rect 315396 488232 315448 488238
rect 315396 488174 315448 488180
rect 313002 487928 313058 487937
rect 313002 487863 313058 487872
rect 313016 487830 313044 487863
rect 312544 487824 312596 487830
rect 312544 487766 312596 487772
rect 313004 487824 313056 487830
rect 313004 487766 313056 487772
rect 312556 487150 312584 487766
rect 319628 487688 319680 487694
rect 319628 487630 319680 487636
rect 318064 487552 318116 487558
rect 318064 487494 318116 487500
rect 318076 487257 318104 487494
rect 319640 487393 319668 487630
rect 320914 487520 320970 487529
rect 322952 487490 322980 488407
rect 326344 487620 326396 487626
rect 326344 487562 326396 487568
rect 324962 487520 325018 487529
rect 320914 487455 320970 487464
rect 322940 487484 322992 487490
rect 319626 487384 319682 487393
rect 320928 487354 320956 487455
rect 324962 487455 325018 487464
rect 322940 487426 322992 487432
rect 319626 487319 319682 487328
rect 320916 487348 320968 487354
rect 318062 487248 318118 487257
rect 318062 487183 318118 487192
rect 319442 487248 319498 487257
rect 319442 487183 319498 487192
rect 299388 487144 299440 487150
rect 299388 487086 299440 487092
rect 311900 487144 311952 487150
rect 311900 487086 311952 487092
rect 312544 487144 312596 487150
rect 312544 487086 312596 487092
rect 311912 464506 311940 487086
rect 318076 472802 318104 487183
rect 318064 472796 318116 472802
rect 318064 472738 318116 472744
rect 311900 464500 311952 464506
rect 311900 464442 311952 464448
rect 319456 460902 319484 487183
rect 319640 479738 319668 487319
rect 320916 487290 320968 487296
rect 320088 487280 320140 487286
rect 320086 487248 320088 487257
rect 320140 487248 320142 487257
rect 320086 487183 320142 487192
rect 320928 485178 320956 487290
rect 322202 487248 322258 487257
rect 321560 487212 321612 487218
rect 322202 487183 322204 487192
rect 321560 487154 321612 487160
rect 322256 487183 322258 487192
rect 322204 487154 322256 487160
rect 320916 485172 320968 485178
rect 320916 485114 320968 485120
rect 321572 482458 321600 487154
rect 322952 486674 322980 487426
rect 324976 487422 325004 487455
rect 324964 487416 325016 487422
rect 324964 487358 325016 487364
rect 324318 487248 324374 487257
rect 324318 487183 324374 487192
rect 322940 486668 322992 486674
rect 322940 486610 322992 486616
rect 321560 482452 321612 482458
rect 321560 482394 321612 482400
rect 319628 479732 319680 479738
rect 319628 479674 319680 479680
rect 324332 472734 324360 487183
rect 324976 474162 325004 487358
rect 326356 487257 326384 487562
rect 326342 487248 326398 487257
rect 326342 487183 326398 487192
rect 329838 487248 329894 487257
rect 329838 487183 329894 487192
rect 335358 487248 335414 487257
rect 335358 487183 335414 487192
rect 339498 487248 339554 487257
rect 339498 487183 339554 487192
rect 345018 487248 345074 487257
rect 345018 487183 345074 487192
rect 349158 487248 349214 487257
rect 349158 487183 349214 487192
rect 354678 487248 354734 487257
rect 354678 487183 354734 487192
rect 360198 487248 360254 487257
rect 360198 487183 360254 487192
rect 326356 476066 326384 487183
rect 326344 476060 326396 476066
rect 326344 476002 326396 476008
rect 329852 475454 329880 487183
rect 329840 475448 329892 475454
rect 329840 475390 329892 475396
rect 324964 474156 325016 474162
rect 324964 474098 325016 474104
rect 335372 474094 335400 487183
rect 339512 479670 339540 487183
rect 339500 479664 339552 479670
rect 339500 479606 339552 479612
rect 335360 474088 335412 474094
rect 335360 474030 335412 474036
rect 324320 472728 324372 472734
rect 324320 472670 324372 472676
rect 345032 463146 345060 487183
rect 345020 463140 345072 463146
rect 345020 463082 345072 463088
rect 349172 461718 349200 487183
rect 354692 478310 354720 487183
rect 360212 482390 360240 487183
rect 360200 482384 360252 482390
rect 360200 482326 360252 482332
rect 354680 478304 354732 478310
rect 354680 478246 354732 478252
rect 395356 478174 395384 699654
rect 395344 478168 395396 478174
rect 395344 478110 395396 478116
rect 399496 468586 399524 700334
rect 403636 476882 403664 700402
rect 405016 489190 405044 700538
rect 429856 700534 429884 703520
rect 409144 700528 409196 700534
rect 409144 700470 409196 700476
rect 429844 700528 429896 700534
rect 429844 700470 429896 700476
rect 406384 700324 406436 700330
rect 406384 700266 406436 700272
rect 405004 489184 405056 489190
rect 405004 489126 405056 489132
rect 403624 476876 403676 476882
rect 403624 476818 403676 476824
rect 399484 468580 399536 468586
rect 399484 468522 399536 468528
rect 406396 465798 406424 700266
rect 407946 636440 408002 636449
rect 407946 636375 408002 636384
rect 407670 635352 407726 635361
rect 407670 635287 407726 635296
rect 407578 628008 407634 628017
rect 407578 627943 407634 627952
rect 407592 598806 407620 627943
rect 407580 598800 407632 598806
rect 407580 598742 407632 598748
rect 406476 596352 406528 596358
rect 406476 596294 406528 596300
rect 406488 478242 406516 596294
rect 407684 585818 407712 635287
rect 407762 632632 407818 632641
rect 407762 632567 407818 632576
rect 407672 585812 407724 585818
rect 407672 585754 407724 585760
rect 407684 526561 407712 585754
rect 407670 526552 407726 526561
rect 407670 526487 407726 526496
rect 407776 523569 407804 632567
rect 407854 607744 407910 607753
rect 407854 607679 407910 607688
rect 407762 523560 407818 523569
rect 407762 523495 407818 523504
rect 407486 521656 407542 521665
rect 407486 521591 407542 521600
rect 407500 520305 407528 521591
rect 407670 520976 407726 520985
rect 407670 520911 407726 520920
rect 407486 520296 407542 520305
rect 407486 520231 407542 520240
rect 407394 517984 407450 517993
rect 407394 517919 407450 517928
rect 407408 488209 407436 517919
rect 407500 488374 407528 520231
rect 407488 488368 407540 488374
rect 407684 488345 407712 520911
rect 407776 489870 407804 523495
rect 407868 498409 407896 607679
rect 407960 598942 407988 636375
rect 408038 633720 408094 633729
rect 408038 633655 408094 633664
rect 408052 600030 408080 633655
rect 408130 631000 408186 631009
rect 408130 630935 408186 630944
rect 408040 600024 408092 600030
rect 408040 599966 408092 599972
rect 407948 598936 408000 598942
rect 407948 598878 408000 598884
rect 408144 598874 408172 630935
rect 408222 629640 408278 629649
rect 408222 629575 408278 629584
rect 408132 598868 408184 598874
rect 408132 598810 408184 598816
rect 408132 596556 408184 596562
rect 408132 596498 408184 596504
rect 408040 596488 408092 596494
rect 408040 596430 408092 596436
rect 407948 596420 408000 596426
rect 407948 596362 408000 596368
rect 407854 498400 407910 498409
rect 407854 498335 407910 498344
rect 407764 489864 407816 489870
rect 407764 489806 407816 489812
rect 407868 488442 407896 498335
rect 407960 488510 407988 596362
rect 407948 488504 408000 488510
rect 407948 488446 408000 488452
rect 407856 488436 407908 488442
rect 407856 488378 407908 488384
rect 407488 488310 407540 488316
rect 407670 488336 407726 488345
rect 407670 488271 407726 488280
rect 407960 488238 407988 488446
rect 408052 488442 408080 596430
rect 408040 488436 408092 488442
rect 408040 488378 408092 488384
rect 408052 488306 408080 488378
rect 408144 488374 408172 596498
rect 408236 521665 408264 629575
rect 408314 610056 408370 610065
rect 408314 609991 408370 610000
rect 408222 521656 408278 521665
rect 408222 521591 408278 521600
rect 408328 500313 408356 609991
rect 408406 608696 408462 608705
rect 408406 608631 408462 608640
rect 408314 500304 408370 500313
rect 408314 500239 408370 500248
rect 408222 498264 408278 498273
rect 408222 498199 408278 498208
rect 408132 488368 408184 488374
rect 408132 488310 408184 488316
rect 408040 488300 408092 488306
rect 408040 488242 408092 488248
rect 407948 488232 408000 488238
rect 407394 488200 407450 488209
rect 407948 488174 408000 488180
rect 407394 488135 407450 488144
rect 408144 487830 408172 488310
rect 408132 487824 408184 487830
rect 408132 487766 408184 487772
rect 406476 478236 406528 478242
rect 406476 478178 406528 478184
rect 406384 465792 406436 465798
rect 406384 465734 406436 465740
rect 408236 463078 408264 498199
rect 408328 488170 408356 500239
rect 408420 498681 408448 608631
rect 408406 498672 408462 498681
rect 408406 498607 408462 498616
rect 408420 498273 408448 498607
rect 408406 498264 408462 498273
rect 408406 498199 408462 498208
rect 408316 488164 408368 488170
rect 408316 488106 408368 488112
rect 409156 467226 409184 700470
rect 462332 700466 462360 703520
rect 462320 700460 462372 700466
rect 462320 700402 462372 700408
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 509884 700324 509936 700330
rect 509884 700266 509936 700272
rect 508504 670744 508556 670750
rect 508504 670686 508556 670692
rect 501604 630692 501656 630698
rect 501604 630634 501656 630640
rect 440238 597544 440294 597553
rect 440238 597479 440294 597488
rect 449898 597544 449954 597553
rect 449898 597479 449954 597488
rect 459558 597544 459614 597553
rect 459558 597479 459614 597488
rect 434718 597408 434774 597417
rect 434718 597343 434774 597352
rect 434732 597310 434760 597343
rect 434720 597304 434772 597310
rect 422574 597272 422630 597281
rect 422574 597207 422630 597216
rect 426438 597272 426494 597281
rect 426438 597207 426494 597216
rect 427818 597272 427874 597281
rect 427818 597207 427820 597216
rect 409418 596864 409474 596873
rect 409418 596799 409474 596808
rect 409328 596284 409380 596290
rect 409328 596226 409380 596232
rect 409236 596216 409288 596222
rect 409236 596158 409288 596164
rect 409248 483750 409276 596158
rect 409340 485110 409368 596226
rect 409432 486538 409460 596799
rect 422588 596562 422616 597207
rect 426452 597174 426480 597207
rect 427872 597207 427874 597216
rect 430578 597272 430634 597281
rect 434720 597246 434772 597252
rect 430578 597207 430634 597216
rect 427820 597178 427872 597184
rect 426440 597168 426492 597174
rect 426440 597110 426492 597116
rect 429198 597136 429254 597145
rect 429198 597071 429200 597080
rect 429252 597071 429254 597080
rect 429200 597042 429252 597048
rect 430592 597038 430620 597207
rect 430580 597032 430632 597038
rect 423678 597000 423734 597009
rect 430580 596974 430632 596980
rect 431958 597000 432014 597009
rect 423678 596935 423734 596944
rect 431958 596935 432014 596944
rect 433338 597000 433394 597009
rect 433338 596935 433394 596944
rect 434718 597000 434774 597009
rect 434718 596935 434720 596944
rect 422576 596556 422628 596562
rect 422576 596498 422628 596504
rect 423692 596494 423720 596935
rect 431972 596902 432000 596935
rect 431960 596896 432012 596902
rect 431960 596838 432012 596844
rect 433352 596834 433380 596935
rect 434772 596935 434774 596944
rect 434720 596906 434772 596912
rect 433340 596828 433392 596834
rect 433340 596770 433392 596776
rect 434718 596728 434774 596737
rect 434718 596663 434774 596672
rect 423680 596488 423732 596494
rect 423680 596430 423732 596436
rect 425058 596456 425114 596465
rect 425058 596391 425060 596400
rect 425112 596391 425114 596400
rect 425060 596362 425112 596368
rect 434732 596358 434760 596663
rect 434720 596352 434772 596358
rect 434720 596294 434772 596300
rect 440252 592686 440280 597479
rect 444378 596728 444434 596737
rect 444378 596663 444434 596672
rect 444392 596290 444420 596663
rect 444380 596284 444432 596290
rect 444380 596226 444432 596232
rect 440240 592680 440292 592686
rect 440240 592622 440292 592628
rect 449912 588606 449940 597479
rect 455418 596320 455474 596329
rect 455418 596255 455474 596264
rect 455432 596222 455460 596255
rect 455420 596216 455472 596222
rect 455420 596158 455472 596164
rect 449900 588600 449952 588606
rect 449900 588542 449952 588548
rect 459572 580310 459600 597479
rect 470598 596320 470654 596329
rect 470598 596255 470654 596264
rect 470612 589937 470640 596255
rect 470598 589928 470654 589937
rect 470598 589863 470654 589872
rect 459560 580304 459612 580310
rect 459560 580246 459612 580252
rect 425060 488504 425112 488510
rect 422574 488472 422630 488481
rect 422574 488407 422630 488416
rect 423678 488472 423734 488481
rect 423678 488407 423680 488416
rect 422588 488374 422616 488407
rect 423732 488407 423734 488416
rect 425058 488472 425060 488481
rect 425112 488472 425114 488481
rect 425058 488407 425114 488416
rect 423680 488378 423732 488384
rect 422576 488368 422628 488374
rect 422576 488310 422628 488316
rect 465078 488336 465134 488345
rect 465078 488271 465134 488280
rect 429198 488200 429254 488209
rect 429198 488135 429254 488144
rect 427818 487792 427874 487801
rect 427818 487727 427874 487736
rect 427832 487694 427860 487727
rect 427820 487688 427872 487694
rect 426438 487656 426494 487665
rect 427820 487630 427872 487636
rect 426438 487591 426494 487600
rect 426452 487558 426480 487591
rect 426440 487552 426492 487558
rect 426440 487494 426492 487500
rect 429212 487286 429240 488135
rect 434718 487656 434774 487665
rect 434718 487591 434720 487600
rect 434772 487591 434774 487600
rect 434720 487562 434772 487568
rect 430578 487520 430634 487529
rect 430578 487455 430634 487464
rect 432142 487520 432198 487529
rect 432142 487455 432198 487464
rect 433338 487520 433394 487529
rect 433338 487455 433340 487464
rect 430592 487354 430620 487455
rect 430580 487348 430632 487354
rect 430580 487290 430632 487296
rect 429200 487280 429252 487286
rect 429200 487222 429252 487228
rect 432156 487218 432184 487455
rect 433392 487455 433394 487464
rect 434718 487520 434774 487529
rect 434718 487455 434774 487464
rect 433340 487426 433392 487432
rect 434732 487422 434760 487455
rect 434720 487416 434772 487422
rect 434720 487358 434772 487364
rect 434718 487248 434774 487257
rect 432144 487212 432196 487218
rect 434718 487183 434774 487192
rect 440238 487248 440294 487257
rect 440238 487183 440294 487192
rect 444378 487248 444434 487257
rect 444378 487183 444434 487192
rect 449898 487248 449954 487257
rect 449898 487183 449954 487192
rect 454682 487248 454738 487257
rect 459558 487248 459614 487257
rect 454682 487183 454738 487192
rect 457444 487212 457496 487218
rect 432144 487154 432196 487160
rect 409420 486532 409472 486538
rect 409420 486474 409472 486480
rect 409328 485104 409380 485110
rect 409328 485046 409380 485052
rect 409236 483744 409288 483750
rect 409236 483686 409288 483692
rect 434732 481030 434760 487183
rect 434720 481024 434772 481030
rect 434720 480966 434772 480972
rect 440252 471306 440280 487183
rect 440240 471300 440292 471306
rect 440240 471242 440292 471248
rect 444392 468518 444420 487183
rect 449912 469946 449940 487183
rect 449900 469940 449952 469946
rect 449900 469882 449952 469888
rect 444380 468512 444432 468518
rect 444380 468454 444432 468460
rect 409144 467220 409196 467226
rect 409144 467162 409196 467168
rect 454696 464438 454724 487183
rect 465092 487218 465120 488271
rect 470598 487248 470654 487257
rect 459558 487183 459614 487192
rect 465080 487212 465132 487218
rect 457444 487154 457496 487160
rect 457456 465730 457484 487154
rect 459572 476814 459600 487183
rect 470598 487183 470654 487192
rect 465080 487154 465132 487160
rect 459560 476808 459612 476814
rect 459560 476750 459612 476756
rect 470612 467158 470640 487183
rect 501616 482322 501644 630634
rect 504364 616888 504416 616894
rect 504364 616830 504416 616836
rect 502984 510672 503036 510678
rect 502984 510614 503036 510620
rect 501604 482316 501656 482322
rect 501604 482258 501656 482264
rect 470600 467152 470652 467158
rect 470600 467094 470652 467100
rect 457444 465724 457496 465730
rect 457444 465666 457496 465672
rect 454684 464432 454736 464438
rect 454684 464374 454736 464380
rect 408224 463072 408276 463078
rect 408224 463014 408276 463020
rect 349160 461712 349212 461718
rect 349160 461654 349212 461660
rect 319444 460896 319496 460902
rect 319444 460838 319496 460844
rect 502996 460222 503024 510614
rect 504376 464370 504404 616830
rect 507124 563100 507176 563106
rect 507124 563042 507176 563048
rect 504364 464364 504416 464370
rect 504364 464306 504416 464312
rect 507136 461650 507164 563042
rect 508516 463010 508544 670686
rect 509896 469878 509924 700266
rect 512644 643136 512696 643142
rect 512644 643078 512696 643084
rect 511264 536852 511316 536858
rect 511264 536794 511316 536800
rect 511276 472666 511304 536794
rect 512656 474026 512684 643078
rect 516784 576904 516836 576910
rect 516784 576846 516836 576852
rect 514024 524476 514076 524482
rect 514024 524418 514076 524424
rect 514036 479534 514064 524418
rect 516796 480962 516824 576846
rect 516784 480956 516836 480962
rect 516784 480898 516836 480904
rect 514024 479528 514076 479534
rect 514024 479470 514076 479476
rect 527192 475386 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 486470 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 542360 486464 542412 486470
rect 542360 486406 542412 486412
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 483682 580304 683839
rect 580264 483676 580316 483682
rect 580264 483618 580316 483624
rect 527180 475380 527232 475386
rect 527180 475322 527232 475328
rect 512644 474020 512696 474026
rect 512644 473962 512696 473968
rect 511264 472660 511316 472666
rect 511264 472602 511316 472608
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 509884 469872 509936 469878
rect 509884 469814 509936 469820
rect 508504 463004 508556 463010
rect 508504 462946 508556 462952
rect 507124 461644 507176 461650
rect 507124 461586 507176 461592
rect 502984 460216 503036 460222
rect 502984 460158 503036 460164
rect 363144 458992 363196 458998
rect 363144 458934 363196 458940
rect 299388 458788 299440 458794
rect 299388 458730 299440 458736
rect 329656 458788 329708 458794
rect 329656 458730 329708 458736
rect 299020 456816 299072 456822
rect 299020 456758 299072 456764
rect 298928 455660 298980 455666
rect 298928 455602 298980 455608
rect 298940 449206 298968 455602
rect 299032 453354 299060 456758
rect 299020 453348 299072 453354
rect 299020 453290 299072 453296
rect 299400 451994 299428 458730
rect 299480 458720 299532 458726
rect 299480 458662 299532 458668
rect 299492 454782 299520 458662
rect 299572 458584 299624 458590
rect 299572 458526 299624 458532
rect 299584 454850 299612 458526
rect 309048 458312 309100 458318
rect 309048 458254 309100 458260
rect 299664 458244 299716 458250
rect 299664 458186 299716 458192
rect 299572 454844 299624 454850
rect 299572 454786 299624 454792
rect 299480 454776 299532 454782
rect 299480 454718 299532 454724
rect 299388 451988 299440 451994
rect 299388 451930 299440 451936
rect 299676 451274 299704 458186
rect 299756 456136 299808 456142
rect 299756 456078 299808 456084
rect 300768 456136 300820 456142
rect 300768 456078 300820 456084
rect 299768 453506 299796 456078
rect 300320 455666 300702 455682
rect 300780 455666 300808 456078
rect 309060 455940 309088 458254
rect 321284 458244 321336 458250
rect 321284 458186 321336 458192
rect 317420 457292 317472 457298
rect 317420 457234 317472 457240
rect 312636 456068 312688 456074
rect 312636 456010 312688 456016
rect 312648 455954 312676 456010
rect 312648 455926 312938 455954
rect 317432 455940 317460 457234
rect 321296 455940 321324 458186
rect 325792 457224 325844 457230
rect 325792 457166 325844 457172
rect 325804 455940 325832 457166
rect 329668 455940 329696 458730
rect 342536 458720 342588 458726
rect 342536 458662 342588 458668
rect 338028 457156 338080 457162
rect 338028 457098 338080 457104
rect 334164 457088 334216 457094
rect 334164 457030 334216 457036
rect 334176 455940 334204 457030
rect 338040 455940 338068 457098
rect 342548 455940 342576 458662
rect 346400 458652 346452 458658
rect 346400 458594 346452 458600
rect 346412 455940 346440 458594
rect 350908 458584 350960 458590
rect 350908 458526 350960 458532
rect 350920 455940 350948 458526
rect 359280 458516 359332 458522
rect 359280 458458 359332 458464
rect 355784 458380 355836 458386
rect 355784 458322 355836 458328
rect 355796 457502 355824 458322
rect 355784 457496 355836 457502
rect 355784 457438 355836 457444
rect 354772 457020 354824 457026
rect 354772 456962 354824 456968
rect 354784 455940 354812 456962
rect 359292 455940 359320 458458
rect 363156 455940 363184 458934
rect 371516 458924 371568 458930
rect 371516 458866 371568 458872
rect 367652 458448 367704 458454
rect 367652 458390 367704 458396
rect 367664 455940 367692 458390
rect 371528 455940 371556 458866
rect 379888 458856 379940 458862
rect 379888 458798 379940 458804
rect 376024 458380 376076 458386
rect 376024 458322 376076 458328
rect 376036 455940 376064 458322
rect 379900 455940 379928 458798
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 383752 456952 383804 456958
rect 383752 456894 383804 456900
rect 383764 455940 383792 456894
rect 385500 456884 385552 456890
rect 385500 456826 385552 456832
rect 385316 456000 385368 456006
rect 385316 455942 385368 455948
rect 385040 455864 385092 455870
rect 385040 455806 385092 455812
rect 384120 455796 384172 455802
rect 384120 455738 384172 455744
rect 300308 455660 300702 455666
rect 300360 455654 300702 455660
rect 300768 455660 300820 455666
rect 300308 455602 300360 455608
rect 300768 455602 300820 455608
rect 384028 455592 384080 455598
rect 304184 455518 304566 455546
rect 384028 455534 384080 455540
rect 304184 455394 304212 455518
rect 299848 455388 299900 455394
rect 299848 455330 299900 455336
rect 304172 455388 304224 455394
rect 304172 455330 304224 455336
rect 299860 454918 299888 455330
rect 299848 454912 299900 454918
rect 299848 454854 299900 454860
rect 383934 454200 383990 454209
rect 383856 454158 383934 454186
rect 299768 453478 299888 453506
rect 299676 451246 299796 451274
rect 299768 450702 299796 451246
rect 299756 450696 299808 450702
rect 299756 450638 299808 450644
rect 298928 449200 298980 449206
rect 298928 449142 298980 449148
rect 299386 448624 299442 448633
rect 299386 448559 299442 448568
rect 298836 446412 298888 446418
rect 298836 446354 298888 446360
rect 299110 446312 299166 446321
rect 299110 446247 299166 446256
rect 298926 446176 298982 446185
rect 298926 446111 298982 446120
rect 298742 446040 298798 446049
rect 298742 445975 298798 445984
rect 298652 398268 298704 398274
rect 298652 398210 298704 398216
rect 296444 365696 296496 365702
rect 296444 365638 296496 365644
rect 296352 259412 296404 259418
rect 296352 259354 296404 259360
rect 296168 219428 296220 219434
rect 296168 219370 296220 219376
rect 298756 113150 298784 445975
rect 298834 443864 298890 443873
rect 298834 443799 298890 443808
rect 298848 193186 298876 443799
rect 298940 233238 298968 446111
rect 299018 443184 299074 443193
rect 299018 443119 299074 443128
rect 298928 233232 298980 233238
rect 298928 233174 298980 233180
rect 299032 206990 299060 443119
rect 299124 325650 299152 446247
rect 299296 444576 299348 444582
rect 299296 444518 299348 444524
rect 299202 443320 299258 443329
rect 299202 443255 299258 443264
rect 299112 325644 299164 325650
rect 299112 325586 299164 325592
rect 299216 273222 299244 443255
rect 299308 379506 299336 444518
rect 299400 398546 299428 448559
rect 299860 446486 299888 453478
rect 299848 446480 299900 446486
rect 299848 446422 299900 446428
rect 299480 445052 299532 445058
rect 299480 444994 299532 445000
rect 299492 422294 299520 444994
rect 299846 442640 299902 442649
rect 299846 442575 299902 442584
rect 299492 422266 299796 422294
rect 299572 401260 299624 401266
rect 299572 401202 299624 401208
rect 299480 401056 299532 401062
rect 299480 400998 299532 401004
rect 299492 400722 299520 400998
rect 299584 400994 299612 401202
rect 299664 401124 299716 401130
rect 299664 401066 299716 401072
rect 299572 400988 299624 400994
rect 299572 400930 299624 400936
rect 299572 400784 299624 400790
rect 299572 400726 299624 400732
rect 299480 400716 299532 400722
rect 299480 400658 299532 400664
rect 299480 399016 299532 399022
rect 299480 398958 299532 398964
rect 299388 398540 299440 398546
rect 299388 398482 299440 398488
rect 299296 379500 299348 379506
rect 299296 379442 299348 379448
rect 299204 273216 299256 273222
rect 299204 273158 299256 273164
rect 299020 206984 299072 206990
rect 299020 206926 299072 206932
rect 298836 193180 298888 193186
rect 298836 193122 298888 193128
rect 298744 113144 298796 113150
rect 298744 113086 298796 113092
rect 296076 100700 296128 100706
rect 296076 100642 296128 100648
rect 298100 83632 298152 83638
rect 298100 83574 298152 83580
rect 296720 20188 296772 20194
rect 296720 20130 296772 20136
rect 296732 16574 296760 20130
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 291396 480 291424 16546
rect 292578 6352 292634 6361
rect 292578 6287 292634 6296
rect 292592 480 292620 6287
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 83574
rect 299492 3482 299520 398958
rect 299584 398682 299612 400726
rect 299676 400654 299704 401066
rect 299664 400648 299716 400654
rect 299664 400590 299716 400596
rect 299768 400466 299796 422266
rect 299860 400790 299888 442575
rect 383856 431954 383884 454158
rect 383934 454135 383990 454144
rect 384040 452305 384068 455534
rect 384026 452296 384082 452305
rect 384026 452231 384082 452240
rect 384132 452146 384160 455738
rect 384212 455728 384264 455734
rect 384212 455670 384264 455676
rect 383948 452118 384160 452146
rect 383948 438705 383976 452118
rect 384224 451274 384252 455670
rect 384304 455524 384356 455530
rect 384304 455466 384356 455472
rect 384040 451246 384252 451274
rect 384040 448225 384068 451246
rect 384026 448216 384082 448225
rect 384026 448151 384082 448160
rect 383934 438696 383990 438705
rect 383934 438631 383990 438640
rect 383856 431926 383976 431954
rect 384316 431934 384344 455466
rect 383948 421705 383976 431926
rect 384304 431928 384356 431934
rect 384304 431870 384356 431876
rect 383934 421696 383990 421705
rect 383934 421631 383990 421640
rect 385052 407561 385080 455806
rect 385224 455660 385276 455666
rect 385224 455602 385276 455608
rect 385130 454064 385186 454073
rect 385130 453999 385186 454008
rect 385144 412321 385172 453999
rect 385236 416401 385264 455602
rect 385328 430001 385356 455942
rect 385408 455932 385460 455938
rect 385408 455874 385460 455880
rect 385420 434081 385448 455874
rect 385512 442921 385540 456826
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580264 455456 580316 455462
rect 580264 455398 580316 455404
rect 385498 442912 385554 442921
rect 385498 442847 385554 442856
rect 385406 434072 385462 434081
rect 385406 434007 385462 434016
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 385314 429992 385370 430001
rect 385314 429927 385370 429936
rect 580276 418305 580304 455398
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 385222 416392 385278 416401
rect 385222 416327 385278 416336
rect 385130 412312 385186 412321
rect 385130 412247 385186 412256
rect 385038 407552 385094 407561
rect 385038 407487 385094 407496
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 385038 403472 385094 403481
rect 385038 403407 385094 403416
rect 299848 400784 299900 400790
rect 299848 400726 299900 400732
rect 307576 400648 307628 400654
rect 311900 400648 311952 400654
rect 307628 400596 307786 400602
rect 307576 400590 307786 400596
rect 324228 400648 324280 400654
rect 313278 400616 313334 400625
rect 311952 400596 312294 400602
rect 311900 400590 312294 400596
rect 307588 400574 307786 400590
rect 311912 400574 312294 400590
rect 340972 400648 341024 400654
rect 332598 400616 332654 400625
rect 324280 400596 324530 400602
rect 324228 400590 324530 400596
rect 324240 400574 324530 400590
rect 313278 400551 313334 400560
rect 332654 400574 332902 400602
rect 382738 400616 382794 400625
rect 341024 400596 341274 400602
rect 340972 400590 341274 400596
rect 340984 400574 341274 400590
rect 332598 400551 332654 400560
rect 382794 400574 383134 400602
rect 382738 400551 382794 400560
rect 299768 400438 300058 400466
rect 303908 398750 303936 400044
rect 303896 398744 303948 398750
rect 303896 398686 303948 398692
rect 299572 398676 299624 398682
rect 299572 398618 299624 398624
rect 310518 396536 310574 396545
rect 310518 396471 310574 396480
rect 305000 394528 305052 394534
rect 305000 394470 305052 394476
rect 299572 391468 299624 391474
rect 299572 391410 299624 391416
rect 299584 3874 299612 391410
rect 300860 351348 300912 351354
rect 300860 351290 300912 351296
rect 300872 16574 300900 351290
rect 303620 18896 303672 18902
rect 303620 18838 303672 18844
rect 303632 16574 303660 18838
rect 305012 16574 305040 394470
rect 307758 86320 307814 86329
rect 307758 86255 307814 86264
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299572 3868 299624 3874
rect 299572 3810 299624 3816
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3810
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303160 7948 303212 7954
rect 303160 7890 303212 7896
rect 303172 480 303200 7890
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 7880 306800 7886
rect 306748 7822 306800 7828
rect 306760 480 306788 7822
rect 307772 3398 307800 86255
rect 307850 19952 307906 19961
rect 307850 19887 307906 19896
rect 307864 16574 307892 19887
rect 310532 16574 310560 396471
rect 311900 25832 311952 25838
rect 311900 25774 311952 25780
rect 311912 16574 311940 25774
rect 313292 16574 313320 400551
rect 383658 400480 383714 400489
rect 383658 400415 383714 400424
rect 316144 398002 316172 400044
rect 320652 398070 320680 400044
rect 329024 398274 329052 400044
rect 331220 398948 331272 398954
rect 331220 398890 331272 398896
rect 329012 398268 329064 398274
rect 329012 398210 329064 398216
rect 320640 398064 320692 398070
rect 320640 398006 320692 398012
rect 316132 397996 316184 398002
rect 316132 397938 316184 397944
rect 324318 397352 324374 397361
rect 324318 397287 324374 397296
rect 322940 394460 322992 394466
rect 322940 394402 322992 394408
rect 316040 389972 316092 389978
rect 316040 389914 316092 389920
rect 314660 20120 314712 20126
rect 314660 20062 314712 20068
rect 307864 16546 307984 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 16546
rect 310242 7576 310298 7585
rect 310242 7511 310298 7520
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 7511
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 20062
rect 316052 16574 316080 389914
rect 317420 352844 317472 352850
rect 317420 352786 317472 352792
rect 317432 16574 317460 352786
rect 321560 352776 321612 352782
rect 321560 352718 321612 352724
rect 318800 25764 318852 25770
rect 318800 25706 318852 25712
rect 318812 16574 318840 25706
rect 321572 16574 321600 352718
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 321572 16546 322152 16574
rect 316236 480 316264 16546
rect 317328 7812 317380 7818
rect 317328 7754 317380 7760
rect 317340 480 317368 7754
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 320916 7744 320968 7750
rect 320916 7686 320968 7692
rect 320928 480 320956 7686
rect 322124 480 322152 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 394402
rect 324332 3398 324360 397287
rect 328458 355328 328514 355337
rect 328458 355263 328514 355272
rect 325698 25664 325754 25673
rect 325698 25599 325754 25608
rect 325712 16574 325740 25599
rect 328472 16574 328500 355263
rect 325712 16546 326384 16574
rect 328472 16546 328776 16574
rect 324412 9308 324464 9314
rect 324412 9250 324464 9256
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 9250
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 327998 9208 328054 9217
rect 327998 9143 328054 9152
rect 328012 480 328040 9143
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 12164 330444 12170
rect 330392 12106 330444 12112
rect 330404 480 330432 12106
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 398890
rect 337396 398857 337424 400044
rect 337382 398848 337438 398857
rect 337382 398783 337438 398792
rect 345768 397934 345796 400044
rect 349632 398342 349660 400044
rect 354140 398721 354168 400044
rect 354126 398712 354182 398721
rect 354126 398647 354182 398656
rect 358004 398410 358032 400044
rect 362512 398478 362540 400044
rect 366376 398614 366404 400044
rect 366364 398608 366416 398614
rect 366364 398550 366416 398556
rect 370884 398546 370912 400044
rect 374748 398682 374776 400044
rect 379256 398818 379284 400044
rect 379244 398812 379296 398818
rect 379244 398754 379296 398760
rect 374736 398676 374788 398682
rect 374736 398618 374788 398624
rect 370872 398540 370924 398546
rect 370872 398482 370924 398488
rect 362500 398472 362552 398478
rect 362500 398414 362552 398420
rect 357992 398404 358044 398410
rect 357992 398346 358044 398352
rect 349620 398336 349672 398342
rect 349620 398278 349672 398284
rect 345756 397928 345808 397934
rect 345756 397870 345808 397876
rect 364338 397216 364394 397225
rect 364338 397151 364394 397160
rect 342260 396908 342312 396914
rect 342260 396850 342312 396856
rect 333980 395684 334032 395690
rect 333980 395626 334032 395632
rect 332600 394392 332652 394398
rect 332600 394334 332652 394340
rect 332612 3398 332640 394334
rect 332692 20052 332744 20058
rect 332692 19994 332744 20000
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 19994
rect 333992 16574 334020 395626
rect 340880 394324 340932 394330
rect 340880 394266 340932 394272
rect 336740 80708 336792 80714
rect 336740 80650 336792 80656
rect 335360 21752 335412 21758
rect 335360 21694 335412 21700
rect 335372 16574 335400 21694
rect 336752 16574 336780 80650
rect 339500 21684 339552 21690
rect 339500 21626 339552 21632
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338672 9240 338724 9246
rect 338672 9182 338724 9188
rect 338684 480 338712 9182
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 21626
rect 340892 16574 340920 394266
rect 342272 16574 342300 396850
rect 347780 394256 347832 394262
rect 347780 394198 347832 394204
rect 343638 84824 343694 84833
rect 343638 84759 343694 84768
rect 343652 16574 343680 84759
rect 346398 21584 346454 21593
rect 346398 21519 346454 21528
rect 346412 16574 346440 21519
rect 347792 16574 347820 394198
rect 357440 389904 357492 389910
rect 357440 389846 357492 389852
rect 353300 354340 353352 354346
rect 353300 354282 353352 354288
rect 349160 21616 349212 21622
rect 349160 21558 349212 21564
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 340984 480 341012 16546
rect 342168 9172 342220 9178
rect 342168 9114 342220 9120
rect 342180 480 342208 9114
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 345754 9072 345810 9081
rect 345754 9007 345810 9016
rect 345768 480 345796 9007
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3398 349200 21558
rect 353312 16574 353340 354282
rect 354680 84856 354732 84862
rect 354680 84798 354732 84804
rect 354692 16574 354720 84798
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 351184 13456 351236 13462
rect 351184 13398 351236 13404
rect 349252 9104 349304 9110
rect 349252 9046 349304 9052
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 9046
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 13398
rect 352840 9036 352892 9042
rect 352840 8978 352892 8984
rect 352852 480 352880 8978
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356336 8968 356388 8974
rect 356336 8910 356388 8916
rect 356348 480 356376 8910
rect 357452 3398 357480 389846
rect 361578 354104 361634 354113
rect 361578 354039 361634 354048
rect 357532 21548 357584 21554
rect 357532 21490 357584 21496
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 21490
rect 360198 21448 360254 21457
rect 360198 21383 360254 21392
rect 360212 16574 360240 21383
rect 361592 16574 361620 354039
rect 364352 16574 364380 397151
rect 365720 394188 365772 394194
rect 365720 394130 365772 394136
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 364352 16546 364656 16574
rect 359464 10668 359516 10674
rect 359464 10610 359516 10616
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 10610
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363510 10568 363566 10577
rect 363510 10503 363566 10512
rect 363524 480 363552 10503
rect 364628 480 364656 16546
rect 365732 3210 365760 394130
rect 382280 394120 382332 394126
rect 382280 394062 382332 394068
rect 365812 391400 365864 391406
rect 365812 391342 365864 391348
rect 365824 3398 365852 391342
rect 367100 352708 367152 352714
rect 367100 352650 367152 352656
rect 367112 16574 367140 352650
rect 379520 352640 379572 352646
rect 379520 352582 379572 352588
rect 372620 177336 372672 177342
rect 372620 177278 372672 177284
rect 371240 21480 371292 21486
rect 371240 21422 371292 21428
rect 367112 16546 367784 16574
rect 365812 3392 365864 3398
rect 365812 3334 365864 3340
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 365732 3182 365852 3210
rect 365824 480 365852 3182
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369400 14816 369452 14822
rect 369400 14758 369452 14764
rect 369412 480 369440 14758
rect 370136 10600 370188 10606
rect 370136 10542 370188 10548
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 10542
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 21422
rect 372632 16574 372660 177278
rect 374000 21412 374052 21418
rect 374000 21354 374052 21360
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3398 374040 21354
rect 378138 21312 378194 21321
rect 378138 21247 378194 21256
rect 378152 16574 378180 21247
rect 378152 16546 378456 16574
rect 376024 16312 376076 16318
rect 376024 16254 376076 16260
rect 374092 10532 374144 10538
rect 374092 10474 374144 10480
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 10474
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16254
rect 377678 10432 377734 10441
rect 377678 10367 377734 10376
rect 377692 480 377720 10367
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 352582
rect 381174 10296 381230 10305
rect 381174 10231 381230 10240
rect 381188 480 381216 10231
rect 382292 3398 382320 394062
rect 382370 22944 382426 22953
rect 382370 22879 382426 22888
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 22879
rect 383672 16574 383700 400415
rect 385052 400110 385080 403407
rect 455418 400344 455474 400353
rect 455418 400279 455474 400288
rect 385040 400104 385092 400110
rect 385040 400046 385092 400052
rect 437480 399152 437532 399158
rect 437480 399094 437532 399100
rect 418802 398440 418858 398449
rect 418802 398375 418858 398384
rect 398838 397080 398894 397089
rect 398838 397015 398894 397024
rect 391940 354272 391992 354278
rect 391940 354214 391992 354220
rect 389180 178696 389232 178702
rect 389180 178638 389232 178644
rect 385040 86352 385092 86358
rect 385040 86294 385092 86300
rect 385052 16574 385080 86294
rect 386420 23112 386472 23118
rect 386420 23054 386472 23060
rect 386432 16574 386460 23054
rect 389192 16574 389220 178638
rect 390560 25696 390612 25702
rect 390560 25638 390612 25644
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 388260 6452 388312 6458
rect 388260 6394 388312 6400
rect 388272 480 388300 6394
rect 389468 480 389496 16546
rect 390572 3210 390600 25638
rect 391952 16574 391980 354214
rect 393320 351280 393372 351286
rect 393320 351222 393372 351228
rect 393332 16574 393360 351222
rect 396080 18828 396132 18834
rect 396080 18770 396132 18776
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 390652 10464 390704 10470
rect 390652 10406 390704 10412
rect 390664 3398 390692 10406
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3334
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395344 10396 395396 10402
rect 395344 10338 395396 10344
rect 395356 480 395384 10338
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 18770
rect 397460 17604 397512 17610
rect 397460 17546 397512 17552
rect 397472 16574 397500 17546
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3398 398880 397015
rect 402980 396840 403032 396846
rect 402980 396782 403032 396788
rect 401600 392828 401652 392834
rect 401600 392770 401652 392776
rect 398930 82104 398986 82113
rect 398930 82039 398986 82048
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 82039
rect 400220 27124 400272 27130
rect 400220 27066 400272 27072
rect 400232 16574 400260 27066
rect 401612 16574 401640 392770
rect 402992 16574 403020 396782
rect 409880 396772 409932 396778
rect 409880 396714 409932 396720
rect 404360 352572 404412 352578
rect 404360 352514 404412 352520
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 352514
rect 407120 27056 407172 27062
rect 407120 26998 407172 27004
rect 406016 12028 406068 12034
rect 406016 11970 406068 11976
rect 406028 480 406056 11970
rect 407132 3398 407160 26998
rect 407212 23044 407264 23050
rect 407212 22986 407264 22992
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 22986
rect 409892 16574 409920 396714
rect 411260 354204 411312 354210
rect 411260 354146 411312 354152
rect 411272 16574 411300 354146
rect 414018 22808 414074 22817
rect 414018 22743 414074 22752
rect 414032 16574 414060 22743
rect 416778 22672 416834 22681
rect 416778 22607 416834 22616
rect 416792 16574 416820 22607
rect 418160 18760 418212 18766
rect 418160 18702 418212 18708
rect 418172 16574 418200 18702
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 414032 16546 414336 16574
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 409144 11960 409196 11966
rect 409144 11902 409196 11908
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 11902
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 412638 11792 412694 11801
rect 412638 11727 412694 11736
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 11727
rect 414308 480 414336 16546
rect 415400 12096 415452 12102
rect 415400 12038 415452 12044
rect 415412 3210 415440 12038
rect 415490 11656 415546 11665
rect 415490 11591 415546 11600
rect 415504 3398 415532 11591
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 3182 415532 3210
rect 415504 480 415532 3182
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3874 418844 398375
rect 431958 396944 432014 396953
rect 431958 396879 432014 396888
rect 423680 351212 423732 351218
rect 423680 351154 423732 351160
rect 422300 83564 422352 83570
rect 422300 83506 422352 83512
rect 420920 83496 420972 83502
rect 420920 83438 420972 83444
rect 420184 11892 420236 11898
rect 420184 11834 420236 11840
rect 418804 3868 418856 3874
rect 418804 3810 418856 3816
rect 420196 480 420224 11834
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 83438
rect 422312 16574 422340 83506
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 423692 1018 423720 351154
rect 429200 334620 429252 334626
rect 429200 334562 429252 334568
rect 427820 87712 427872 87718
rect 427820 87654 427872 87660
rect 425060 25628 425112 25634
rect 425060 25570 425112 25576
rect 425072 16574 425100 25570
rect 427832 16574 427860 87654
rect 425072 16546 425744 16574
rect 427832 16546 428504 16574
rect 423772 11824 423824 11830
rect 423772 11766 423824 11772
rect 423680 1012 423732 1018
rect 423680 954 423732 960
rect 423784 480 423812 11766
rect 424968 1012 425020 1018
rect 424968 954 425020 960
rect 424980 480 425008 954
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426808 11756 426860 11762
rect 426808 11698 426860 11704
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 11698
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 334562
rect 430856 13388 430908 13394
rect 430856 13330 430908 13336
rect 430868 480 430896 13330
rect 431972 1170 432000 396879
rect 434718 352880 434774 352889
rect 434718 352815 434774 352824
rect 432050 24440 432106 24449
rect 432050 24375 432106 24384
rect 432064 3398 432092 24375
rect 434732 16574 434760 352815
rect 436100 305652 436152 305658
rect 436100 305594 436152 305600
rect 436112 16574 436140 305594
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433982 13152 434038 13161
rect 433982 13087 434038 13096
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 13087
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 399094
rect 452658 396808 452714 396817
rect 452658 396743 452714 396752
rect 440240 394052 440292 394058
rect 440240 393994 440292 394000
rect 438860 389836 438912 389842
rect 438860 389778 438912 389784
rect 438872 16574 438900 389778
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 393994
rect 445760 354136 445812 354142
rect 445760 354078 445812 354084
rect 443000 186992 443052 186998
rect 443000 186934 443052 186940
rect 441620 22976 441672 22982
rect 441620 22918 441672 22924
rect 441632 16574 441660 22918
rect 443012 16574 443040 186934
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 440332 13320 440384 13326
rect 440332 13262 440384 13268
rect 440344 3398 440372 13262
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445024 13252 445076 13258
rect 445024 13194 445076 13200
rect 445036 480 445064 13194
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 354078
rect 449900 336048 449952 336054
rect 449900 335990 449952 335996
rect 447140 26988 447192 26994
rect 447140 26930 447192 26936
rect 447152 16574 447180 26930
rect 448520 22908 448572 22914
rect 448520 22850 448572 22856
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 1018 448560 22850
rect 449912 16574 449940 335990
rect 452672 16574 452700 396743
rect 454040 86284 454092 86290
rect 454040 86226 454092 86232
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 448612 13184 448664 13190
rect 448612 13126 448664 13132
rect 448520 1012 448572 1018
rect 448520 954 448572 960
rect 448624 480 448652 13126
rect 449808 1012 449860 1018
rect 449808 954 449860 960
rect 449820 480 449848 954
rect 450924 480 450952 16546
rect 451646 13016 451702 13025
rect 451646 12951 451702 12960
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 12951
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 86226
rect 455432 16574 455460 400279
rect 580000 400178 580028 404903
rect 579988 400172 580040 400178
rect 579988 400114 580040 400120
rect 494058 398304 494114 398313
rect 494058 398239 494114 398248
rect 492680 393984 492732 393990
rect 492680 393926 492732 393932
rect 483020 392760 483072 392766
rect 483020 392702 483072 392708
rect 460940 188352 460992 188358
rect 460940 188294 460992 188300
rect 456800 29640 456852 29646
rect 456800 29582 456852 29588
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 29582
rect 456892 22840 456944 22846
rect 456892 22782 456944 22788
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 22782
rect 459560 22772 459612 22778
rect 459560 22714 459612 22720
rect 459572 16574 459600 22714
rect 460952 16574 460980 188294
rect 474740 31068 474792 31074
rect 474740 31010 474792 31016
rect 471980 26920 472032 26926
rect 471980 26862 472032 26868
rect 463700 24472 463752 24478
rect 463700 24414 463752 24420
rect 463712 16574 463740 24414
rect 466458 24304 466514 24313
rect 466458 24239 466514 24248
rect 466472 16574 466500 24239
rect 470598 24168 470654 24177
rect 470598 24103 470654 24112
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 459192 13116 459244 13122
rect 459192 13058 459244 13064
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 13058
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 462320 14748 462372 14754
rect 462320 14690 462372 14696
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 14690
rect 463988 480 464016 16546
rect 465816 14680 465868 14686
rect 465816 14622 465868 14628
rect 465172 3800 465224 3806
rect 465172 3742 465224 3748
rect 465184 480 465212 3742
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 14622
rect 467484 480 467512 16546
rect 469862 14784 469918 14793
rect 469862 14719 469918 14728
rect 468668 3732 468720 3738
rect 468668 3674 468720 3680
rect 468680 480 468708 3674
rect 469876 480 469904 14719
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 24103
rect 471992 16574 472020 26862
rect 473360 24404 473412 24410
rect 473360 24346 473412 24352
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3602 473400 24346
rect 474752 16574 474780 31010
rect 477500 24336 477552 24342
rect 477500 24278 477552 24284
rect 477512 16574 477540 24278
rect 481640 24268 481692 24274
rect 481640 24210 481692 24216
rect 474752 16546 475792 16574
rect 477512 16546 478184 16574
rect 473452 14612 473504 14618
rect 473452 14554 473504 14560
rect 473360 3596 473412 3602
rect 473360 3538 473412 3544
rect 473464 480 473492 14554
rect 474188 3596 474240 3602
rect 474188 3538 474240 3544
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3538
rect 475764 480 475792 16546
rect 476488 14544 476540 14550
rect 476488 14486 476540 14492
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 14486
rect 478156 480 478184 16546
rect 479340 3732 479392 3738
rect 479340 3674 479392 3680
rect 479352 480 479380 3674
rect 480536 3664 480588 3670
rect 480536 3606 480588 3612
rect 480548 480 480576 3606
rect 481652 3602 481680 24210
rect 483032 16574 483060 392702
rect 485778 352744 485834 352753
rect 485778 352679 485834 352688
rect 485792 16574 485820 352679
rect 487158 26888 487214 26897
rect 487158 26823 487214 26832
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 481732 14476 481784 14482
rect 481732 14418 481784 14424
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 14418
rect 482468 3596 482520 3602
rect 482468 3538 482520 3544
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3538
rect 484044 480 484072 16546
rect 484766 14648 484822 14657
rect 484766 14583 484822 14592
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 14583
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 26823
rect 490012 24200 490064 24206
rect 490012 24142 490064 24148
rect 488814 14512 488870 14521
rect 488814 14447 488870 14456
rect 488828 480 488856 14447
rect 490024 6914 490052 24142
rect 492692 16574 492720 393926
rect 494072 16574 494100 398239
rect 543740 398200 543792 398206
rect 507858 398168 507914 398177
rect 543740 398142 543792 398148
rect 507858 398103 507914 398112
rect 498200 392692 498252 392698
rect 498200 392634 498252 392640
rect 496820 24132 496872 24138
rect 496820 24074 496872 24080
rect 496832 16574 496860 24074
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 492312 7676 492364 7682
rect 492312 7618 492364 7624
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3528 491168 3534
rect 491116 3470 491168 3476
rect 491128 480 491156 3470
rect 492324 480 492352 7618
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 495440 16244 495492 16250
rect 495440 16186 495492 16192
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 16186
rect 497108 480 497136 16546
rect 498212 480 498240 392634
rect 506480 355496 506532 355502
rect 506480 355438 506532 355444
rect 503718 86184 503774 86193
rect 503718 86119 503774 86128
rect 499580 82136 499632 82142
rect 499580 82078 499632 82084
rect 499592 16574 499620 82078
rect 499592 16546 500632 16574
rect 498936 16176 498988 16182
rect 498936 16118 498988 16124
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16118
rect 500604 480 500632 16546
rect 502984 16108 503036 16114
rect 502984 16050 503036 16056
rect 501788 3460 501840 3466
rect 501788 3402 501840 3408
rect 501800 480 501828 3402
rect 502996 480 503024 16050
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 86119
rect 506492 3534 506520 355438
rect 506570 352608 506626 352617
rect 506570 352543 506626 352552
rect 506480 3528 506532 3534
rect 505374 3496 505430 3505
rect 506480 3470 506532 3476
rect 505374 3431 505430 3440
rect 505388 480 505416 3431
rect 506584 3346 506612 352543
rect 507872 16574 507900 398103
rect 525798 398032 525854 398041
rect 525798 397967 525854 397976
rect 521658 396672 521714 396681
rect 521658 396607 521714 396616
rect 512000 392624 512052 392630
rect 512000 392566 512052 392572
rect 510620 355428 510672 355434
rect 510620 355370 510672 355376
rect 510632 16574 510660 355370
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 509608 16040 509660 16046
rect 509608 15982 509660 15988
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 15982
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 392566
rect 514760 391332 514812 391338
rect 514760 391274 514812 391280
rect 513380 15972 513432 15978
rect 513380 15914 513432 15920
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 15914
rect 514772 3534 514800 391274
rect 514852 356856 514904 356862
rect 514852 356798 514904 356804
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 356798
rect 517520 356788 517572 356794
rect 517520 356730 517572 356736
rect 517532 16574 517560 356730
rect 517532 16546 517928 16574
rect 517152 15904 517204 15910
rect 517152 15846 517204 15852
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 15846
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 520278 16008 520334 16017
rect 520278 15943 520334 15952
rect 519544 5160 519596 5166
rect 519544 5102 519596 5108
rect 519556 480 519584 5102
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 15943
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 396607
rect 525812 16574 525840 397967
rect 535460 395616 535512 395622
rect 535460 395558 535512 395564
rect 529940 391264 529992 391270
rect 529940 391206 529992 391212
rect 527180 17536 527232 17542
rect 527180 17478 527232 17484
rect 527192 16574 527220 17478
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523774 15872 523830 15881
rect 523774 15807 523830 15816
rect 523038 5128 523094 5137
rect 523038 5063 523094 5072
rect 523052 480 523080 5063
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 15807
rect 525432 5092 525484 5098
rect 525432 5034 525484 5040
rect 525444 480 525472 5034
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 529020 7608 529072 7614
rect 529020 7550 529072 7556
rect 529032 480 529060 7550
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 529952 354 529980 391206
rect 531320 356720 531372 356726
rect 531320 356662 531372 356668
rect 531332 3534 531360 356662
rect 531412 87644 531464 87650
rect 531412 87586 531464 87592
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 87586
rect 534080 17468 534132 17474
rect 534080 17410 534132 17416
rect 534092 16574 534120 17410
rect 535472 16574 535500 395558
rect 542360 354068 542412 354074
rect 542360 354010 542412 354016
rect 538218 353968 538274 353977
rect 538218 353903 538274 353912
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 533712 5024 533764 5030
rect 533712 4966 533764 4972
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 4966
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 537220 480 537248 4898
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 353903
rect 540978 17504 541034 17513
rect 540978 17439 541034 17448
rect 540992 16574 541020 17439
rect 542372 16574 542400 354010
rect 543752 16574 543780 398142
rect 564440 398132 564492 398138
rect 564440 398074 564492 398080
rect 549260 395548 549312 395554
rect 549260 395490 549312 395496
rect 546500 354000 546552 354006
rect 546500 353942 546552 353948
rect 545120 17400 545172 17406
rect 545120 17342 545172 17348
rect 545132 16574 545160 17342
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 539598 8936 539654 8945
rect 539598 8871 539654 8880
rect 539612 480 539640 8871
rect 540794 4992 540850 5001
rect 540794 4927 540850 4936
rect 540808 480 540836 4927
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 353942
rect 547880 17332 547932 17338
rect 547880 17274 547932 17280
rect 547892 16574 547920 17274
rect 549272 16574 549300 395490
rect 560300 395480 560352 395486
rect 560300 395422 560352 395428
rect 556158 395312 556214 395321
rect 556158 395247 556214 395256
rect 550640 355360 550692 355366
rect 550640 355302 550692 355308
rect 550652 16574 550680 355302
rect 552020 17264 552072 17270
rect 552020 17206 552072 17212
rect 552032 16574 552060 17206
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 547880 4888 547932 4894
rect 547880 4830 547932 4836
rect 547892 480 547920 4830
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553768 10328 553820 10334
rect 553768 10270 553820 10276
rect 553780 480 553808 10270
rect 554964 4820 555016 4826
rect 554964 4762 555016 4768
rect 554976 480 555004 4762
rect 556172 3534 556200 395247
rect 556250 17368 556306 17377
rect 556250 17303 556306 17312
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 17303
rect 558918 17232 558974 17241
rect 558918 17167 558974 17176
rect 558932 16574 558960 17167
rect 560312 16574 560340 395422
rect 563060 18692 563112 18698
rect 563060 18634 563112 18640
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 558550 4856 558606 4865
rect 558550 4791 558606 4800
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 4791
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562048 6384 562100 6390
rect 562048 6326 562100 6332
rect 562060 480 562088 6326
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 18634
rect 564452 3534 564480 398074
rect 564532 395412 564584 395418
rect 564532 395354 564584 395360
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 395354
rect 571340 395344 571392 395350
rect 571340 395286 571392 395292
rect 567200 25560 567252 25566
rect 567200 25502 567252 25508
rect 567212 16574 567240 25502
rect 569960 18624 570012 18630
rect 569960 18566 570012 18572
rect 569972 16574 570000 18566
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 566832 6316 566884 6322
rect 566832 6258 566884 6264
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 6258
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 6248 569184 6254
rect 569132 6190 569184 6196
rect 569144 480 569172 6190
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 395286
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 572720 348424 572772 348430
rect 572720 348366 572772 348372
rect 572732 16574 572760 348366
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 582380 191140 582432 191146
rect 582380 191082 582432 191088
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 581092 167680 581144 167686
rect 581092 167622 581144 167628
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 576858 87544 576914 87553
rect 576858 87479 576914 87488
rect 574098 25528 574154 25537
rect 574098 25463 574154 25472
rect 574112 16574 574140 25463
rect 576872 16574 576900 87479
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 578240 19984 578292 19990
rect 578240 19926 578292 19932
rect 578252 16574 578280 19926
rect 581104 16574 581132 167622
rect 582392 16574 582420 191082
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 572720 6180 572772 6186
rect 572720 6122 572772 6128
rect 572732 480 572760 6122
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576306 6216 576362 6225
rect 576306 6151 576362 6160
rect 576320 480 576348 6151
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 581000 3868 581052 3874
rect 581000 3810 581052 3816
rect 579802 3360 579858 3369
rect 579802 3295 579858 3304
rect 579816 480 579844 3295
rect 581012 480 581040 3810
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 566888 3386 566944
rect 3146 553832 3202 553888
rect 3330 527856 3386 527912
rect 3238 501744 3294 501800
rect 3238 475632 3294 475688
rect 2870 462576 2926 462632
rect 3238 449520 3294 449576
rect 3514 671200 3570 671256
rect 3606 658144 3662 658200
rect 3698 632032 3754 632088
rect 3790 619112 3846 619168
rect 3882 606056 3938 606112
rect 3974 579944 4030 580000
rect 4066 514800 4122 514856
rect 78586 636384 78642 636440
rect 78310 635296 78366 635352
rect 78218 633664 78274 633720
rect 77758 632576 77814 632632
rect 78126 630944 78182 631000
rect 77850 629584 77906 629640
rect 77758 523504 77814 523560
rect 78034 627952 78090 628008
rect 77942 608640 77998 608696
rect 77850 520240 77906 520296
rect 78402 610000 78458 610056
rect 78494 607688 78550 607744
rect 102874 597488 102930 597544
rect 106186 597488 106242 597544
rect 92478 597352 92534 597408
rect 99286 597352 99342 597408
rect 102046 597352 102102 597408
rect 94042 596944 94098 597000
rect 97906 596964 97962 597000
rect 97906 596944 97908 596964
rect 97908 596944 97960 596964
rect 97960 596944 97962 596964
rect 78494 526632 78550 526688
rect 78310 526496 78366 526552
rect 78310 523640 78366 523696
rect 78126 520920 78182 520976
rect 78034 499840 78090 499896
rect 77942 498616 77998 498672
rect 78402 498344 78458 498400
rect 78586 517928 78642 517984
rect 100666 597080 100722 597136
rect 103426 597216 103482 597272
rect 106094 597236 106150 597272
rect 106094 597216 106096 597236
rect 106096 597216 106148 597236
rect 106148 597216 106150 597236
rect 104806 597100 104862 597136
rect 104806 597080 104808 597100
rect 104808 597080 104860 597100
rect 104860 597080 104862 597100
rect 95238 596264 95294 596320
rect 131026 596944 131082 597000
rect 126886 596672 126942 596728
rect 136546 596536 136602 596592
rect 140686 596556 140742 596592
rect 140686 596536 140688 596556
rect 140688 596536 140740 596556
rect 140740 596536 140742 596556
rect 115846 596264 115902 596320
rect 121366 596284 121422 596320
rect 121366 596264 121368 596284
rect 121368 596264 121420 596284
rect 121420 596264 121422 596284
rect 92938 488452 92940 488472
rect 92940 488452 92992 488472
rect 92992 488452 92994 488472
rect 92938 488416 92994 488452
rect 94226 488436 94282 488472
rect 94226 488416 94228 488436
rect 94228 488416 94280 488436
rect 94280 488416 94282 488436
rect 95330 488416 95386 488472
rect 97814 488416 97870 488472
rect 98918 488416 98974 488472
rect 100022 488416 100078 488472
rect 101126 488416 101182 488472
rect 102414 488416 102470 488472
rect 104806 488416 104862 488472
rect 105726 488416 105782 488472
rect 103426 488008 103482 488064
rect 106002 488144 106058 488200
rect 111706 488144 111762 488200
rect 115846 487192 115902 487248
rect 121366 487192 121422 487248
rect 126886 487192 126942 487248
rect 131026 487192 131082 487248
rect 136546 487192 136602 487248
rect 140686 487192 140742 487248
rect 173254 596808 173310 596864
rect 3146 423580 3148 423600
rect 3148 423580 3200 423600
rect 3200 423580 3202 423600
rect 3146 423544 3202 423580
rect 3238 410488 3294 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 319232 3386 319288
rect 2778 306212 2780 306232
rect 2780 306212 2832 306232
rect 2832 306212 2834 306232
rect 2778 306176 2834 306212
rect 3146 267144 3202 267200
rect 3054 214920 3110 214976
rect 2778 201864 2834 201920
rect 3054 162832 3110 162888
rect 2778 149776 2834 149832
rect 3330 110608 3386 110664
rect 2778 97552 2834 97608
rect 3330 71576 3386 71632
rect 4066 345344 4122 345400
rect 3974 293120 4030 293176
rect 3882 241032 3938 241088
rect 3790 188808 3846 188864
rect 3698 136720 3754 136776
rect 3606 84632 3662 84688
rect 3514 58520 3570 58576
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 187330 637064 187386 637120
rect 186778 635976 186834 636032
rect 186686 630264 186742 630320
rect 186870 634344 186926 634400
rect 187238 631624 187294 631680
rect 187146 628632 187202 628688
rect 187054 610272 187110 610328
rect 186962 608368 187018 608424
rect 186778 525952 186834 526008
rect 186870 524320 186926 524376
rect 186686 520240 186742 520296
rect 186778 517520 186834 517576
rect 187422 633256 187478 633312
rect 187330 527040 187386 527096
rect 187606 608640 187662 608696
rect 187514 524320 187570 524376
rect 187422 523232 187478 523288
rect 187238 521600 187294 521656
rect 187146 518608 187202 518664
rect 187146 517520 187202 517576
rect 187054 500248 187110 500304
rect 186962 498344 187018 498400
rect 188434 525952 188490 526008
rect 187606 498616 187662 498672
rect 207110 597488 207166 597544
rect 208398 597488 208454 597544
rect 210054 597488 210110 597544
rect 211158 597488 211214 597544
rect 212446 597488 212502 597544
rect 213826 597488 213882 597544
rect 214838 597488 214894 597544
rect 215298 597488 215354 597544
rect 215942 597488 215998 597544
rect 226246 597488 226302 597544
rect 235906 597488 235962 597544
rect 245566 597488 245622 597544
rect 251086 597488 251142 597544
rect 204350 597080 204406 597136
rect 202878 596400 202934 596456
rect 204258 596264 204314 596320
rect 219438 596264 219494 596320
rect 189078 498616 189134 498672
rect 231766 597216 231822 597272
rect 241426 596808 241482 596864
rect 204442 488436 204498 488472
rect 204442 488416 204444 488436
rect 204444 488416 204496 488436
rect 204496 488416 204498 488436
rect 214838 488416 214894 488472
rect 202878 488180 202880 488200
rect 202880 488180 202932 488200
rect 202932 488180 202934 488200
rect 202878 488144 202934 488180
rect 211158 488280 211214 488336
rect 213734 488280 213790 488336
rect 215390 488280 215446 488336
rect 211802 487464 211858 487520
rect 210422 487348 210478 487384
rect 210422 487328 210424 487348
rect 210424 487328 210476 487348
rect 210476 487328 210478 487348
rect 203522 487192 203578 487248
rect 204902 487192 204958 487248
rect 207662 487212 207718 487248
rect 207662 487192 207664 487212
rect 207664 487192 207716 487212
rect 207716 487192 207718 487212
rect 209042 487228 209044 487248
rect 209044 487228 209096 487248
rect 209096 487228 209098 487248
rect 209042 487192 209098 487228
rect 216586 487192 216642 487248
rect 213182 446256 213238 446312
rect 11058 396616 11114 396672
rect 570 8880 626 8936
rect 13818 177248 13874 177304
rect 25502 397976 25558 398032
rect 13542 14456 13598 14512
rect 17038 11600 17094 11656
rect 64878 396752 64934 396808
rect 27710 395256 27766 395312
rect 28998 392536 29054 392592
rect 45558 395392 45614 395448
rect 49698 177384 49754 177440
rect 48502 12960 48558 13016
rect 51354 9016 51410 9072
rect 63498 177520 63554 177576
rect 67638 395528 67694 395584
rect 66718 13096 66774 13152
rect 84198 15816 84254 15872
rect 81622 14592 81678 14648
rect 83278 10240 83334 10296
rect 86406 10376 86462 10432
rect 178682 398248 178738 398304
rect 102138 355272 102194 355328
rect 100758 10512 100814 10568
rect 118698 395664 118754 395720
rect 120078 177656 120134 177712
rect 118790 11736 118846 11792
rect 122286 11872 122342 11928
rect 139398 393896 139454 393952
rect 138846 15952 138902 16008
rect 137650 6160 137706 6216
rect 151818 396888 151874 396944
rect 153198 352552 153254 352608
rect 155222 14728 155278 14784
rect 175278 351056 175334 351112
rect 170770 7520 170826 7576
rect 174266 7656 174322 7712
rect 173162 6296 173218 6352
rect 188342 398112 188398 398168
rect 187698 392672 187754 392728
rect 192022 7792 192078 7848
rect 190826 6432 190882 6488
rect 212078 446120 212134 446176
rect 210422 445984 210478 446040
rect 210238 445032 210294 445088
rect 209686 444896 209742 444952
rect 209502 444352 209558 444408
rect 210054 444624 210110 444680
rect 209962 443944 210018 444000
rect 210606 444488 210662 444544
rect 211710 444080 211766 444136
rect 211618 443808 211674 443864
rect 211250 443672 211306 443728
rect 209410 443536 209466 443592
rect 212262 444080 212318 444136
rect 212814 444080 212870 444136
rect 211986 443400 212042 443456
rect 220726 487192 220782 487248
rect 220082 443944 220138 444000
rect 212722 443400 212778 443456
rect 215850 443420 215906 443456
rect 215850 443400 215852 443420
rect 215852 443400 215904 443420
rect 215904 443400 215906 443420
rect 216586 443420 216642 443456
rect 226246 487192 226302 487248
rect 224406 448568 224462 448624
rect 225694 454008 225750 454064
rect 227166 446528 227222 446584
rect 226246 445848 226302 445904
rect 231766 487192 231822 487248
rect 229190 446800 229246 446856
rect 229006 446664 229062 446720
rect 229742 446392 229798 446448
rect 216586 443400 216588 443420
rect 216588 443400 216640 443420
rect 216640 443400 216642 443420
rect 220082 443400 220138 443456
rect 230386 446528 230442 446584
rect 231398 445032 231454 445088
rect 232134 454280 232190 454336
rect 235906 487192 235962 487248
rect 241426 487192 241482 487248
rect 244646 487192 244702 487248
rect 232686 454144 232742 454200
rect 234066 449792 234122 449848
rect 234250 449656 234306 449712
rect 234526 449656 234582 449712
rect 249982 487192 250038 487248
rect 250902 444080 250958 444136
rect 255410 449520 255466 449576
rect 255502 446392 255558 446448
rect 256422 449520 256478 449576
rect 256606 446548 256662 446584
rect 256606 446528 256608 446548
rect 256608 446528 256660 446548
rect 256660 446528 256662 446548
rect 264978 446664 265034 446720
rect 256422 444080 256478 444136
rect 256790 445712 256846 445768
rect 207754 398792 207810 398848
rect 202142 398384 202198 398440
rect 194414 6568 194470 6624
rect 203614 397704 203670 397760
rect 206190 7928 206246 7984
rect 208398 392808 208454 392864
rect 210330 397432 210386 397488
rect 210330 397024 210386 397080
rect 210330 396752 210386 396808
rect 210698 397976 210754 398032
rect 210698 397704 210754 397760
rect 211158 398248 211214 398304
rect 211526 398520 211582 398576
rect 211434 397568 211490 397624
rect 211618 397704 211674 397760
rect 211342 397432 211398 397488
rect 211250 396752 211306 396808
rect 211894 397840 211950 397896
rect 211802 397568 211858 397624
rect 212170 398248 212226 398304
rect 212262 397840 212318 397896
rect 212446 398248 212502 398304
rect 212538 397704 212594 397760
rect 212630 397432 212686 397488
rect 212814 397976 212870 398032
rect 212998 397568 213054 397624
rect 213366 398384 213422 398440
rect 213274 394712 213330 394768
rect 214010 398792 214066 398848
rect 214194 397704 214250 397760
rect 214286 397568 214342 397624
rect 214102 397432 214158 397488
rect 213918 395392 213974 395448
rect 215298 397432 215354 397488
rect 215574 397704 215630 397760
rect 215482 397568 215538 397624
rect 215390 397024 215446 397080
rect 215850 397840 215906 397896
rect 215942 393760 215998 393816
rect 215758 393488 215814 393544
rect 216678 397568 216734 397624
rect 216954 398656 217010 398712
rect 217046 397840 217102 397896
rect 216862 397704 216918 397760
rect 216770 397432 216826 397488
rect 217230 398792 217286 398848
rect 217506 398792 217562 398848
rect 217690 398792 217746 398848
rect 218058 397568 218114 397624
rect 218242 397704 218298 397760
rect 218150 397432 218206 397488
rect 219346 399064 219402 399120
rect 219346 398656 219402 398712
rect 219530 397432 219586 397488
rect 219806 397568 219862 397624
rect 219714 397432 219770 397488
rect 219622 395664 219678 395720
rect 220910 397704 220966 397760
rect 221002 397568 221058 397624
rect 221186 397568 221242 397624
rect 221094 397432 221150 397488
rect 222198 397704 222254 397760
rect 222290 397432 222346 397488
rect 223578 397704 223634 397760
rect 223854 397568 223910 397624
rect 223762 397432 223818 397488
rect 223946 397432 224002 397488
rect 224958 397840 225014 397896
rect 225142 397568 225198 397624
rect 225418 397704 225474 397760
rect 225234 397432 225290 397488
rect 226522 397568 226578 397624
rect 226338 397432 226394 397488
rect 229006 397568 229062 397624
rect 228914 397432 228970 397488
rect 229374 398928 229430 398984
rect 229190 398112 229246 398168
rect 229742 398112 229798 398168
rect 230202 397840 230258 397896
rect 230110 397568 230166 397624
rect 230386 397704 230442 397760
rect 230294 397432 230350 397488
rect 231582 397704 231638 397760
rect 231766 397568 231822 397624
rect 231674 397432 231730 397488
rect 232134 396480 232190 396536
rect 232594 396752 232650 396808
rect 232962 397840 233018 397896
rect 232870 397568 232926 397624
rect 233146 397704 233202 397760
rect 233054 397432 233110 397488
rect 234434 397704 234490 397760
rect 234342 397568 234398 397624
rect 234250 397432 234306 397488
rect 234710 399880 234766 399936
rect 234434 396480 234490 396536
rect 235722 397568 235778 397624
rect 235906 397704 235962 397760
rect 235814 397432 235870 397488
rect 235630 397296 235686 397352
rect 237102 397704 237158 397760
rect 237286 397568 237342 397624
rect 237194 397432 237250 397488
rect 238574 397704 238630 397760
rect 238482 397568 238538 397624
rect 238390 397432 238446 397488
rect 238666 397160 238722 397216
rect 238850 396752 238906 396808
rect 239126 396752 239182 396808
rect 239770 397568 239826 397624
rect 239678 397432 239734 397488
rect 240046 397704 240102 397760
rect 239954 397432 240010 397488
rect 240230 399880 240286 399936
rect 241334 397432 241390 397488
rect 241426 397024 241482 397080
rect 242622 398112 242678 398168
rect 242530 397704 242586 397760
rect 242438 397568 242494 397624
rect 237378 5344 237434 5400
rect 239310 3712 239366 3768
rect 240506 3576 240562 3632
rect 242806 397840 242862 397896
rect 242714 397432 242770 397488
rect 244002 397568 244058 397624
rect 244186 397704 244242 397760
rect 243910 396888 243966 396944
rect 244094 397432 244150 397488
rect 245382 398928 245438 398984
rect 245474 397432 245530 397488
rect 245750 399880 245806 399936
rect 245566 396752 245622 396808
rect 246210 398248 246266 398304
rect 246486 398656 246542 398712
rect 246762 397840 246818 397896
rect 246670 397568 246726 397624
rect 246946 397704 247002 397760
rect 246854 397432 246910 397488
rect 247038 397024 247094 397080
rect 247038 396616 247094 396672
rect 247314 398520 247370 398576
rect 247314 398248 247370 398304
rect 247958 398248 248014 398304
rect 248142 397840 248198 397896
rect 248234 397704 248290 397760
rect 248326 397568 248382 397624
rect 248050 397432 248106 397488
rect 248510 398656 248566 398712
rect 248510 398384 248566 398440
rect 248786 398248 248842 398304
rect 248786 398112 248842 398168
rect 242898 3440 242954 3496
rect 249062 398384 249118 398440
rect 249522 397568 249578 397624
rect 249706 397704 249762 397760
rect 249614 397432 249670 397488
rect 249890 398112 249946 398168
rect 250810 397568 250866 397624
rect 251086 397704 251142 397760
rect 250994 397432 251050 397488
rect 250902 396616 250958 396672
rect 251270 397976 251326 398032
rect 252190 397704 252246 397760
rect 252282 397568 252338 397624
rect 252466 397840 252522 397896
rect 252374 397432 252430 397488
rect 253662 399200 253718 399256
rect 253570 397568 253626 397624
rect 253846 397704 253902 397760
rect 253754 397432 253810 397488
rect 255042 397568 255098 397624
rect 255226 397704 255282 397760
rect 255134 397432 255190 397488
rect 255226 395392 255282 395448
rect 255410 398384 255466 398440
rect 255962 398656 256018 398712
rect 254674 5208 254730 5264
rect 257342 395528 257398 395584
rect 260102 397840 260158 397896
rect 291934 449520 291990 449576
rect 265806 444896 265862 444952
rect 265622 444760 265678 444816
rect 265714 443400 265770 443456
rect 265898 443672 265954 443728
rect 257066 3304 257122 3360
rect 271142 398520 271198 398576
rect 273258 177248 273314 177304
rect 274822 6432 274878 6488
rect 276110 18536 276166 18592
rect 283562 444624 283618 444680
rect 292946 442720 293002 442776
rect 293130 400968 293186 401024
rect 292946 400832 293002 400888
rect 293406 488008 293462 488064
rect 297914 636928 297970 636984
rect 297822 634208 297878 634264
rect 297638 633120 297694 633176
rect 297454 631488 297510 631544
rect 296994 610136 297050 610192
rect 296902 608232 296958 608288
rect 296810 521464 296866 521520
rect 297086 608640 297142 608696
rect 296994 500792 297050 500848
rect 297178 525952 297234 526008
rect 297086 498616 297142 498672
rect 296902 498208 296958 498264
rect 296810 488280 296866 488336
rect 297546 628496 297602 628552
rect 297362 524320 297418 524376
rect 297270 521600 297326 521656
rect 297270 520240 297326 520296
rect 297454 521464 297510 521520
rect 297730 630128 297786 630184
rect 297638 523232 297694 523288
rect 297546 518608 297602 518664
rect 297546 517520 297602 517576
rect 297362 489776 297418 489832
rect 298006 635840 298062 635896
rect 318338 597488 318394 597544
rect 319442 597488 319498 597544
rect 320086 597488 320142 597544
rect 320914 597488 320970 597544
rect 322294 597488 322350 597544
rect 322938 597488 322994 597544
rect 324318 597488 324374 597544
rect 325790 597488 325846 597544
rect 329838 597488 329894 597544
rect 345018 597488 345074 597544
rect 360198 597488 360254 597544
rect 314658 596944 314714 597000
rect 313278 596828 313334 596864
rect 313278 596808 313280 596828
rect 313280 596808 313332 596828
rect 313332 596808 313334 596828
rect 298006 527060 298062 527096
rect 298006 527040 298008 527060
rect 298008 527040 298060 527060
rect 298060 527040 298062 527060
rect 297730 521600 297786 521656
rect 298006 517520 298062 517576
rect 297914 500792 297970 500848
rect 297914 500248 297970 500304
rect 297822 498208 297878 498264
rect 298006 488144 298062 488200
rect 297362 449792 297418 449848
rect 297178 449656 297234 449712
rect 296074 444488 296130 444544
rect 295982 442312 296038 442368
rect 291198 393896 291254 393952
rect 289818 20168 289874 20224
rect 292578 20032 292634 20088
rect 296166 442176 296222 442232
rect 296350 442448 296406 442504
rect 297822 452376 297878 452432
rect 298006 448296 298062 448352
rect 298098 446392 298154 446448
rect 297178 434696 297234 434752
rect 298006 443536 298062 443592
rect 298006 439456 298062 439512
rect 298006 430616 298062 430672
rect 298006 425856 298062 425912
rect 297546 421776 297602 421832
rect 297454 417016 297510 417072
rect 297362 412936 297418 412992
rect 298006 408176 298062 408232
rect 298006 404096 298062 404152
rect 311898 596536 311954 596592
rect 324410 597352 324466 597408
rect 339498 596944 339554 597000
rect 335358 596264 335414 596320
rect 349158 597080 349214 597136
rect 354678 596264 354734 596320
rect 314290 488416 314346 488472
rect 315394 488416 315450 488472
rect 322938 488416 322994 488472
rect 313002 487872 313058 487928
rect 320914 487464 320970 487520
rect 319626 487328 319682 487384
rect 324962 487464 325018 487520
rect 318062 487192 318118 487248
rect 319442 487192 319498 487248
rect 320086 487228 320088 487248
rect 320088 487228 320140 487248
rect 320140 487228 320142 487248
rect 320086 487192 320142 487228
rect 322202 487212 322258 487248
rect 322202 487192 322204 487212
rect 322204 487192 322256 487212
rect 322256 487192 322258 487212
rect 324318 487192 324374 487248
rect 326342 487192 326398 487248
rect 329838 487192 329894 487248
rect 335358 487192 335414 487248
rect 339498 487192 339554 487248
rect 345018 487192 345074 487248
rect 349158 487192 349214 487248
rect 354678 487192 354734 487248
rect 360198 487192 360254 487248
rect 407946 636384 408002 636440
rect 407670 635296 407726 635352
rect 407578 627952 407634 628008
rect 407762 632576 407818 632632
rect 407670 526496 407726 526552
rect 407854 607688 407910 607744
rect 407762 523504 407818 523560
rect 407486 521600 407542 521656
rect 407670 520920 407726 520976
rect 407486 520240 407542 520296
rect 407394 517928 407450 517984
rect 408038 633664 408094 633720
rect 408130 630944 408186 631000
rect 408222 629584 408278 629640
rect 407854 498344 407910 498400
rect 407670 488280 407726 488336
rect 408314 610000 408370 610056
rect 408222 521600 408278 521656
rect 408406 608640 408462 608696
rect 408314 500248 408370 500304
rect 408222 498208 408278 498264
rect 407394 488144 407450 488200
rect 408406 498616 408462 498672
rect 408406 498208 408462 498264
rect 440238 597488 440294 597544
rect 449898 597488 449954 597544
rect 459558 597488 459614 597544
rect 434718 597352 434774 597408
rect 422574 597216 422630 597272
rect 426438 597216 426494 597272
rect 427818 597236 427874 597272
rect 427818 597216 427820 597236
rect 427820 597216 427872 597236
rect 427872 597216 427874 597236
rect 409418 596808 409474 596864
rect 430578 597216 430634 597272
rect 429198 597100 429254 597136
rect 429198 597080 429200 597100
rect 429200 597080 429252 597100
rect 429252 597080 429254 597100
rect 423678 596944 423734 597000
rect 431958 596944 432014 597000
rect 433338 596944 433394 597000
rect 434718 596964 434774 597000
rect 434718 596944 434720 596964
rect 434720 596944 434772 596964
rect 434772 596944 434774 596964
rect 434718 596672 434774 596728
rect 425058 596420 425114 596456
rect 425058 596400 425060 596420
rect 425060 596400 425112 596420
rect 425112 596400 425114 596420
rect 444378 596672 444434 596728
rect 455418 596264 455474 596320
rect 470598 596264 470654 596320
rect 470598 589872 470654 589928
rect 422574 488416 422630 488472
rect 423678 488436 423734 488472
rect 423678 488416 423680 488436
rect 423680 488416 423732 488436
rect 423732 488416 423734 488436
rect 425058 488452 425060 488472
rect 425060 488452 425112 488472
rect 425112 488452 425114 488472
rect 425058 488416 425114 488452
rect 465078 488280 465134 488336
rect 429198 488144 429254 488200
rect 427818 487736 427874 487792
rect 426438 487600 426494 487656
rect 434718 487620 434774 487656
rect 434718 487600 434720 487620
rect 434720 487600 434772 487620
rect 434772 487600 434774 487620
rect 430578 487464 430634 487520
rect 432142 487464 432198 487520
rect 433338 487484 433394 487520
rect 433338 487464 433340 487484
rect 433340 487464 433392 487484
rect 433392 487464 433394 487484
rect 434718 487464 434774 487520
rect 434718 487192 434774 487248
rect 440238 487192 440294 487248
rect 444378 487192 444434 487248
rect 449898 487192 449954 487248
rect 454682 487192 454738 487248
rect 459558 487192 459614 487248
rect 470598 487192 470654 487248
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 299386 448568 299442 448624
rect 299110 446256 299166 446312
rect 298926 446120 298982 446176
rect 298742 445984 298798 446040
rect 298834 443808 298890 443864
rect 299018 443128 299074 443184
rect 299202 443264 299258 443320
rect 299846 442584 299902 442640
rect 292578 6296 292634 6352
rect 383934 454144 383990 454200
rect 384026 452240 384082 452296
rect 384026 448160 384082 448216
rect 383934 438640 383990 438696
rect 383934 421640 383990 421696
rect 385130 454008 385186 454064
rect 385498 442856 385554 442912
rect 385406 434016 385462 434072
rect 580170 431568 580226 431624
rect 385314 429936 385370 429992
rect 580262 418240 580318 418296
rect 385222 416336 385278 416392
rect 385130 412256 385186 412312
rect 385038 407496 385094 407552
rect 579986 404912 580042 404968
rect 385038 403416 385094 403472
rect 313278 400560 313334 400616
rect 332598 400560 332654 400616
rect 382738 400560 382794 400616
rect 310518 396480 310574 396536
rect 307758 86264 307814 86320
rect 307850 19896 307906 19952
rect 383658 400424 383714 400480
rect 324318 397296 324374 397352
rect 310242 7520 310298 7576
rect 328458 355272 328514 355328
rect 325698 25608 325754 25664
rect 327998 9152 328054 9208
rect 337382 398792 337438 398848
rect 354126 398656 354182 398712
rect 364338 397160 364394 397216
rect 343638 84768 343694 84824
rect 346398 21528 346454 21584
rect 345754 9016 345810 9072
rect 361578 354048 361634 354104
rect 360198 21392 360254 21448
rect 363510 10512 363566 10568
rect 378138 21256 378194 21312
rect 377678 10376 377734 10432
rect 381174 10240 381230 10296
rect 382370 22888 382426 22944
rect 455418 400288 455474 400344
rect 418802 398384 418858 398440
rect 398838 397024 398894 397080
rect 398930 82048 398986 82104
rect 414018 22752 414074 22808
rect 416778 22616 416834 22672
rect 412638 11736 412694 11792
rect 415490 11600 415546 11656
rect 431958 396888 432014 396944
rect 434718 352824 434774 352880
rect 432050 24384 432106 24440
rect 433982 13096 434038 13152
rect 452658 396752 452714 396808
rect 451646 12960 451702 13016
rect 494058 398248 494114 398304
rect 466458 24248 466514 24304
rect 470598 24112 470654 24168
rect 469862 14728 469918 14784
rect 485778 352688 485834 352744
rect 487158 26832 487214 26888
rect 484766 14592 484822 14648
rect 488814 14456 488870 14512
rect 507858 398112 507914 398168
rect 503718 86128 503774 86184
rect 506570 352552 506626 352608
rect 505374 3440 505430 3496
rect 525798 397976 525854 398032
rect 521658 396616 521714 396672
rect 520278 15952 520334 16008
rect 523774 15816 523830 15872
rect 523038 5072 523094 5128
rect 538218 353912 538274 353968
rect 540978 17448 541034 17504
rect 539598 8880 539654 8936
rect 540794 4936 540850 4992
rect 556158 395256 556214 395312
rect 556250 17312 556306 17368
rect 558918 17176 558974 17232
rect 558550 4800 558606 4856
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 576858 87488 576914 87544
rect 574098 25472 574154 25528
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 576306 6160 576362 6216
rect 579802 3304 579858 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3601 658202 3667 658205
rect -960 658200 3667 658202
rect -960 658144 3606 658200
rect 3662 658144 3667 658200
rect -960 658142 3667 658144
rect -960 658052 480 658142
rect 3601 658139 3667 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 187325 637122 187391 637125
rect 187325 637120 189458 637122
rect 187325 637064 187330 637120
rect 187386 637064 189458 637120
rect 187325 637062 189458 637064
rect 187325 637059 187391 637062
rect 189398 637060 189458 637062
rect 78581 636442 78647 636445
rect 80002 636442 80062 637030
rect 189398 637000 190072 637060
rect 299430 637000 300012 637060
rect 297909 636986 297975 636989
rect 299430 636986 299490 637000
rect 297909 636984 299490 636986
rect 297909 636928 297914 636984
rect 297970 636928 299490 636984
rect 297909 636926 299490 636928
rect 297909 636923 297975 636926
rect 78581 636440 80062 636442
rect 78581 636384 78586 636440
rect 78642 636384 80062 636440
rect 78581 636382 80062 636384
rect 407941 636442 408007 636445
rect 410002 636442 410062 637030
rect 407941 636440 410062 636442
rect 407941 636384 407946 636440
rect 408002 636384 410062 636440
rect 407941 636382 410062 636384
rect 78581 636379 78647 636382
rect 407941 636379 408007 636382
rect 186773 636034 186839 636037
rect 186773 636032 189458 636034
rect 186773 635976 186778 636032
rect 186834 635976 189458 636032
rect 186773 635974 189458 635976
rect 186773 635971 186839 635974
rect 189398 635972 189458 635974
rect 78305 635354 78371 635357
rect 80002 635354 80062 635942
rect 189398 635912 190072 635972
rect 299430 635912 300012 635972
rect 298001 635898 298067 635901
rect 299430 635898 299490 635912
rect 298001 635896 299490 635898
rect 298001 635840 298006 635896
rect 298062 635840 299490 635896
rect 298001 635838 299490 635840
rect 298001 635835 298067 635838
rect 78305 635352 80062 635354
rect 78305 635296 78310 635352
rect 78366 635296 80062 635352
rect 78305 635294 80062 635296
rect 407665 635354 407731 635357
rect 410002 635354 410062 635942
rect 407665 635352 410062 635354
rect 407665 635296 407670 635352
rect 407726 635296 410062 635352
rect 407665 635294 410062 635296
rect 78305 635291 78371 635294
rect 407665 635291 407731 635294
rect 186865 634402 186931 634405
rect 186865 634400 189458 634402
rect 186865 634344 186870 634400
rect 186926 634344 189458 634400
rect 186865 634342 189458 634344
rect 186865 634339 186931 634342
rect 189398 634340 189458 634342
rect 78213 633722 78279 633725
rect 80002 633722 80062 634310
rect 189398 634280 190072 634340
rect 299430 634280 300012 634340
rect 297817 634266 297883 634269
rect 299430 634266 299490 634280
rect 297817 634264 299490 634266
rect 297817 634208 297822 634264
rect 297878 634208 299490 634264
rect 297817 634206 299490 634208
rect 297817 634203 297883 634206
rect 78213 633720 80062 633722
rect 78213 633664 78218 633720
rect 78274 633664 80062 633720
rect 78213 633662 80062 633664
rect 408033 633722 408099 633725
rect 410002 633722 410062 634310
rect 408033 633720 410062 633722
rect 408033 633664 408038 633720
rect 408094 633664 410062 633720
rect 408033 633662 410062 633664
rect 78213 633659 78279 633662
rect 408033 633659 408099 633662
rect 187417 633314 187483 633317
rect 187417 633312 189458 633314
rect 187417 633256 187422 633312
rect 187478 633256 189458 633312
rect 187417 633254 189458 633256
rect 187417 633251 187483 633254
rect 189398 633252 189458 633254
rect 77753 632634 77819 632637
rect 80002 632634 80062 633222
rect 189398 633192 190072 633252
rect 299430 633192 300012 633252
rect 297633 633178 297699 633181
rect 299430 633178 299490 633192
rect 297633 633176 299490 633178
rect 297633 633120 297638 633176
rect 297694 633120 299490 633176
rect 297633 633118 299490 633120
rect 297633 633115 297699 633118
rect 77753 632632 80062 632634
rect 77753 632576 77758 632632
rect 77814 632576 80062 632632
rect 77753 632574 80062 632576
rect 407757 632634 407823 632637
rect 410002 632634 410062 633222
rect 407757 632632 410062 632634
rect 407757 632576 407762 632632
rect 407818 632576 410062 632632
rect 407757 632574 410062 632576
rect 77753 632571 77819 632574
rect 407757 632571 407823 632574
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 187233 631682 187299 631685
rect 187233 631680 189458 631682
rect 187233 631624 187238 631680
rect 187294 631624 189458 631680
rect 187233 631622 189458 631624
rect 187233 631619 187299 631622
rect 189398 631620 189458 631622
rect 78121 631002 78187 631005
rect 80002 631002 80062 631590
rect 189398 631560 190072 631620
rect 299430 631560 300012 631620
rect 297449 631546 297515 631549
rect 299430 631546 299490 631560
rect 297449 631544 299490 631546
rect 297449 631488 297454 631544
rect 297510 631488 299490 631544
rect 297449 631486 299490 631488
rect 297449 631483 297515 631486
rect 78121 631000 80062 631002
rect 78121 630944 78126 631000
rect 78182 630944 80062 631000
rect 78121 630942 80062 630944
rect 408125 631002 408191 631005
rect 410002 631002 410062 631590
rect 408125 631000 410062 631002
rect 408125 630944 408130 631000
rect 408186 630944 410062 631000
rect 408125 630942 410062 630944
rect 78121 630939 78187 630942
rect 408125 630939 408191 630942
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect 186681 630322 186747 630325
rect 186681 630320 189458 630322
rect 186681 630264 186686 630320
rect 186742 630264 189458 630320
rect 186681 630262 189458 630264
rect 186681 630259 186747 630262
rect 189398 630260 189458 630262
rect 77845 629642 77911 629645
rect 80002 629642 80062 630230
rect 189398 630200 190072 630260
rect 299430 630200 300012 630260
rect 297725 630186 297791 630189
rect 299430 630186 299490 630200
rect 297725 630184 299490 630186
rect 297725 630128 297730 630184
rect 297786 630128 299490 630184
rect 297725 630126 299490 630128
rect 297725 630123 297791 630126
rect 77845 629640 80062 629642
rect 77845 629584 77850 629640
rect 77906 629584 80062 629640
rect 77845 629582 80062 629584
rect 408217 629642 408283 629645
rect 410002 629642 410062 630230
rect 408217 629640 410062 629642
rect 408217 629584 408222 629640
rect 408278 629584 410062 629640
rect 408217 629582 410062 629584
rect 77845 629579 77911 629582
rect 408217 629579 408283 629582
rect 187141 628690 187207 628693
rect 187141 628688 189458 628690
rect 187141 628632 187146 628688
rect 187202 628632 189458 628688
rect 187141 628630 189458 628632
rect 187141 628627 187207 628630
rect 189398 628628 189458 628630
rect 78029 628010 78095 628013
rect 80002 628010 80062 628598
rect 189398 628568 190072 628628
rect 299430 628568 300012 628628
rect 297541 628554 297607 628557
rect 299430 628554 299490 628568
rect 297541 628552 299490 628554
rect 297541 628496 297546 628552
rect 297602 628496 299490 628552
rect 297541 628494 299490 628496
rect 297541 628491 297607 628494
rect 78029 628008 80062 628010
rect 78029 627952 78034 628008
rect 78090 627952 80062 628008
rect 78029 627950 80062 627952
rect 407573 628010 407639 628013
rect 410002 628010 410062 628598
rect 407573 628008 410062 628010
rect 407573 627952 407578 628008
rect 407634 627952 410062 628008
rect 407573 627950 410062 627952
rect 78029 627947 78095 627950
rect 407573 627947 407639 627950
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 187049 610330 187115 610333
rect 187049 610328 189458 610330
rect 187049 610272 187054 610328
rect 187110 610272 189458 610328
rect 187049 610270 189458 610272
rect 187049 610267 187115 610270
rect 189398 610268 189458 610270
rect 78397 610058 78463 610061
rect 80002 610058 80062 610238
rect 189398 610208 190072 610268
rect 299430 610208 300012 610268
rect 296989 610194 297055 610197
rect 299430 610194 299490 610208
rect 296989 610192 299490 610194
rect 296989 610136 296994 610192
rect 297050 610136 299490 610192
rect 296989 610134 299490 610136
rect 296989 610131 297055 610134
rect 78397 610056 80062 610058
rect 78397 610000 78402 610056
rect 78458 610000 80062 610056
rect 78397 609998 80062 610000
rect 408309 610058 408375 610061
rect 410002 610058 410062 610238
rect 408309 610056 410062 610058
rect 408309 610000 408314 610056
rect 408370 610000 410062 610056
rect 408309 609998 410062 610000
rect 78397 609995 78463 609998
rect 408309 609995 408375 609998
rect 77937 608698 78003 608701
rect 187601 608698 187667 608701
rect 297081 608698 297147 608701
rect 408401 608698 408467 608701
rect 77937 608696 80062 608698
rect 77937 608640 77942 608696
rect 77998 608640 80062 608696
rect 77937 608638 80062 608640
rect 77937 608635 78003 608638
rect 80002 608606 80062 608638
rect 187601 608696 189458 608698
rect 187601 608640 187606 608696
rect 187662 608640 189458 608696
rect 187601 608638 189458 608640
rect 187601 608635 187667 608638
rect 189398 608636 189458 608638
rect 297081 608696 299490 608698
rect 297081 608640 297086 608696
rect 297142 608640 299490 608696
rect 297081 608638 299490 608640
rect 189398 608576 190072 608636
rect 297081 608635 297147 608638
rect 299430 608636 299490 608638
rect 408401 608696 410062 608698
rect 408401 608640 408406 608696
rect 408462 608640 410062 608696
rect 408401 608638 410062 608640
rect 299430 608576 300012 608636
rect 408401 608635 408467 608638
rect 410002 608606 410062 608638
rect 186957 608426 187023 608429
rect 186957 608424 189458 608426
rect 186957 608368 186962 608424
rect 187018 608368 189458 608424
rect 186957 608366 189458 608368
rect 186957 608363 187023 608366
rect 189398 608364 189458 608366
rect 78489 607746 78555 607749
rect 80002 607746 80062 608334
rect 189398 608304 190072 608364
rect 299430 608304 300012 608364
rect 296897 608290 296963 608293
rect 299430 608290 299490 608304
rect 296897 608288 299490 608290
rect 296897 608232 296902 608288
rect 296958 608232 299490 608288
rect 296897 608230 299490 608232
rect 296897 608227 296963 608230
rect 78489 607744 80062 607746
rect 78489 607688 78494 607744
rect 78550 607688 80062 607744
rect 78489 607686 80062 607688
rect 407849 607746 407915 607749
rect 410002 607746 410062 608334
rect 407849 607744 410062 607746
rect 407849 607688 407854 607744
rect 407910 607688 410062 607744
rect 407849 607686 410062 607688
rect 78489 607683 78555 607686
rect 407849 607683 407915 607686
rect -960 606114 480 606204
rect 3877 606114 3943 606117
rect -960 606112 3943 606114
rect -960 606056 3882 606112
rect 3938 606056 3943 606112
rect -960 606054 3943 606056
rect -960 605964 480 606054
rect 3877 606051 3943 606054
rect 583520 604060 584960 604300
rect 102358 597484 102364 597548
rect 102428 597546 102434 597548
rect 102869 597546 102935 597549
rect 102428 597544 102935 597546
rect 102428 597488 102874 597544
rect 102930 597488 102935 597544
rect 102428 597486 102935 597488
rect 102428 597484 102434 597486
rect 102869 597483 102935 597486
rect 105302 597484 105308 597548
rect 105372 597546 105378 597548
rect 106181 597546 106247 597549
rect 105372 597544 106247 597546
rect 105372 597488 106186 597544
rect 106242 597488 106247 597544
rect 105372 597486 106247 597488
rect 105372 597484 105378 597486
rect 106181 597483 106247 597486
rect 207105 597546 207171 597549
rect 207606 597546 207612 597548
rect 207105 597544 207612 597546
rect 207105 597488 207110 597544
rect 207166 597488 207612 597544
rect 207105 597486 207612 597488
rect 207105 597483 207171 597486
rect 207606 597484 207612 597486
rect 207676 597484 207682 597548
rect 208393 597546 208459 597549
rect 210049 597548 210115 597549
rect 211153 597548 211219 597549
rect 212441 597548 212507 597549
rect 208894 597546 208900 597548
rect 208393 597544 208900 597546
rect 208393 597488 208398 597544
rect 208454 597488 208900 597544
rect 208393 597486 208900 597488
rect 208393 597483 208459 597486
rect 208894 597484 208900 597486
rect 208964 597484 208970 597548
rect 209998 597546 210004 597548
rect 209958 597486 210004 597546
rect 210068 597544 210115 597548
rect 211102 597546 211108 597548
rect 210110 597488 210115 597544
rect 209998 597484 210004 597486
rect 210068 597484 210115 597488
rect 211062 597486 211108 597546
rect 211172 597544 211219 597548
rect 212390 597546 212396 597548
rect 211214 597488 211219 597544
rect 211102 597484 211108 597486
rect 211172 597484 211219 597488
rect 212350 597486 212396 597546
rect 212460 597544 212507 597548
rect 212502 597488 212507 597544
rect 212390 597484 212396 597486
rect 212460 597484 212507 597488
rect 213494 597484 213500 597548
rect 213564 597546 213570 597548
rect 213821 597546 213887 597549
rect 214833 597548 214899 597549
rect 214782 597546 214788 597548
rect 213564 597544 213887 597546
rect 213564 597488 213826 597544
rect 213882 597488 213887 597544
rect 213564 597486 213887 597488
rect 214742 597486 214788 597546
rect 214852 597544 214899 597548
rect 215293 597548 215359 597549
rect 215293 597546 215340 597548
rect 214894 597488 214899 597544
rect 213564 597484 213570 597486
rect 210049 597483 210115 597484
rect 211153 597483 211219 597484
rect 212441 597483 212507 597484
rect 213821 597483 213887 597486
rect 214782 597484 214788 597486
rect 214852 597484 214899 597488
rect 215248 597544 215340 597546
rect 215248 597488 215298 597544
rect 215248 597486 215340 597488
rect 214833 597483 214899 597484
rect 215293 597484 215340 597486
rect 215404 597484 215410 597548
rect 215702 597484 215708 597548
rect 215772 597546 215778 597548
rect 215937 597546 216003 597549
rect 215772 597544 216003 597546
rect 215772 597488 215942 597544
rect 215998 597488 216003 597544
rect 215772 597486 216003 597488
rect 215772 597484 215778 597486
rect 215293 597483 215359 597484
rect 215937 597483 216003 597486
rect 225454 597484 225460 597548
rect 225524 597546 225530 597548
rect 226241 597546 226307 597549
rect 225524 597544 226307 597546
rect 225524 597488 226246 597544
rect 226302 597488 226307 597544
rect 225524 597486 226307 597488
rect 225524 597484 225530 597486
rect 226241 597483 226307 597486
rect 235574 597484 235580 597548
rect 235644 597546 235650 597548
rect 235901 597546 235967 597549
rect 245561 597548 245627 597549
rect 235644 597544 235967 597546
rect 235644 597488 235906 597544
rect 235962 597488 235967 597544
rect 235644 597486 235967 597488
rect 235644 597484 235650 597486
rect 235901 597483 235967 597486
rect 245510 597484 245516 597548
rect 245580 597546 245627 597548
rect 245580 597544 245672 597546
rect 245622 597488 245672 597544
rect 245580 597486 245672 597488
rect 245580 597484 245627 597486
rect 250478 597484 250484 597548
rect 250548 597546 250554 597548
rect 251081 597546 251147 597549
rect 250548 597544 251147 597546
rect 250548 597488 251086 597544
rect 251142 597488 251147 597544
rect 250548 597486 251147 597488
rect 250548 597484 250554 597486
rect 245561 597483 245627 597484
rect 251081 597483 251147 597486
rect 317638 597484 317644 597548
rect 317708 597546 317714 597548
rect 318333 597546 318399 597549
rect 317708 597544 318399 597546
rect 317708 597488 318338 597544
rect 318394 597488 318399 597544
rect 317708 597486 318399 597488
rect 317708 597484 317714 597486
rect 318333 597483 318399 597486
rect 318926 597484 318932 597548
rect 318996 597546 319002 597548
rect 319437 597546 319503 597549
rect 320081 597548 320147 597549
rect 320030 597546 320036 597548
rect 318996 597544 319503 597546
rect 318996 597488 319442 597544
rect 319498 597488 319503 597544
rect 318996 597486 319503 597488
rect 319990 597486 320036 597546
rect 320100 597544 320147 597548
rect 320142 597488 320147 597544
rect 318996 597484 319002 597486
rect 319437 597483 319503 597486
rect 320030 597484 320036 597486
rect 320100 597484 320147 597488
rect 320081 597483 320147 597484
rect 320909 597546 320975 597549
rect 322289 597548 322355 597549
rect 321134 597546 321140 597548
rect 320909 597544 321140 597546
rect 320909 597488 320914 597544
rect 320970 597488 321140 597544
rect 320909 597486 321140 597488
rect 320909 597483 320975 597486
rect 321134 597484 321140 597486
rect 321204 597484 321210 597548
rect 322238 597546 322244 597548
rect 322198 597486 322244 597546
rect 322308 597544 322355 597548
rect 322350 597488 322355 597544
rect 322238 597484 322244 597486
rect 322308 597484 322355 597488
rect 322289 597483 322355 597484
rect 322933 597546 322999 597549
rect 323342 597546 323348 597548
rect 322933 597544 323348 597546
rect 322933 597488 322938 597544
rect 322994 597488 323348 597544
rect 322933 597486 323348 597488
rect 322933 597483 322999 597486
rect 323342 597484 323348 597486
rect 323412 597484 323418 597548
rect 324313 597546 324379 597549
rect 325785 597548 325851 597549
rect 325182 597546 325188 597548
rect 324313 597544 325188 597546
rect 324313 597488 324318 597544
rect 324374 597488 325188 597544
rect 324313 597486 325188 597488
rect 324313 597483 324379 597486
rect 325182 597484 325188 597486
rect 325252 597484 325258 597548
rect 325734 597546 325740 597548
rect 325694 597486 325740 597546
rect 325804 597544 325851 597548
rect 325846 597488 325851 597544
rect 325734 597484 325740 597486
rect 325804 597484 325851 597488
rect 325785 597483 325851 597484
rect 329833 597546 329899 597549
rect 330518 597546 330524 597548
rect 329833 597544 330524 597546
rect 329833 597488 329838 597544
rect 329894 597488 330524 597544
rect 329833 597486 330524 597488
rect 329833 597483 329899 597486
rect 330518 597484 330524 597486
rect 330588 597484 330594 597548
rect 345013 597546 345079 597549
rect 345606 597546 345612 597548
rect 345013 597544 345612 597546
rect 345013 597488 345018 597544
rect 345074 597488 345612 597544
rect 345013 597486 345612 597488
rect 345013 597483 345079 597486
rect 345606 597484 345612 597486
rect 345676 597484 345682 597548
rect 360193 597546 360259 597549
rect 360510 597546 360516 597548
rect 360193 597544 360516 597546
rect 360193 597488 360198 597544
rect 360254 597488 360516 597544
rect 360193 597486 360516 597488
rect 360193 597483 360259 597486
rect 360510 597484 360516 597486
rect 360580 597484 360586 597548
rect 440233 597546 440299 597549
rect 440366 597546 440372 597548
rect 440233 597544 440372 597546
rect 440233 597488 440238 597544
rect 440294 597488 440372 597544
rect 440233 597486 440372 597488
rect 440233 597483 440299 597486
rect 440366 597484 440372 597486
rect 440436 597484 440442 597548
rect 449893 597546 449959 597549
rect 450486 597546 450492 597548
rect 449893 597544 450492 597546
rect 449893 597488 449898 597544
rect 449954 597488 450492 597544
rect 449893 597486 450492 597488
rect 449893 597483 449959 597486
rect 450486 597484 450492 597486
rect 450556 597484 450562 597548
rect 459553 597546 459619 597549
rect 460422 597546 460428 597548
rect 459553 597544 460428 597546
rect 459553 597488 459558 597544
rect 459614 597488 460428 597544
rect 459553 597486 460428 597488
rect 459553 597483 459619 597486
rect 460422 597484 460428 597486
rect 460492 597484 460498 597548
rect 92473 597410 92539 597413
rect 92974 597410 92980 597412
rect 92473 597408 92980 597410
rect 92473 597352 92478 597408
rect 92534 597352 92980 597408
rect 92473 597350 92980 597352
rect 92473 597347 92539 597350
rect 92974 597348 92980 597350
rect 93044 597348 93050 597412
rect 98862 597348 98868 597412
rect 98932 597410 98938 597412
rect 99281 597410 99347 597413
rect 98932 597408 99347 597410
rect 98932 597352 99286 597408
rect 99342 597352 99347 597408
rect 98932 597350 99347 597352
rect 98932 597348 98938 597350
rect 99281 597347 99347 597350
rect 101070 597348 101076 597412
rect 101140 597410 101146 597412
rect 102041 597410 102107 597413
rect 101140 597408 102107 597410
rect 101140 597352 102046 597408
rect 102102 597352 102107 597408
rect 101140 597350 102107 597352
rect 101140 597348 101146 597350
rect 102041 597347 102107 597350
rect 324405 597410 324471 597413
rect 324814 597410 324820 597412
rect 324405 597408 324820 597410
rect 324405 597352 324410 597408
rect 324466 597352 324820 597408
rect 324405 597350 324820 597352
rect 324405 597347 324471 597350
rect 324814 597348 324820 597350
rect 324884 597348 324890 597412
rect 434713 597410 434779 597413
rect 435582 597410 435588 597412
rect 434713 597408 435588 597410
rect 434713 597352 434718 597408
rect 434774 597352 435588 597408
rect 434713 597350 435588 597352
rect 434713 597347 434779 597350
rect 435582 597348 435588 597350
rect 435652 597348 435658 597412
rect 103278 597212 103284 597276
rect 103348 597274 103354 597276
rect 103421 597274 103487 597277
rect 103348 597272 103487 597274
rect 103348 597216 103426 597272
rect 103482 597216 103487 597272
rect 103348 597214 103487 597216
rect 103348 597212 103354 597214
rect 103421 597211 103487 597214
rect 105670 597212 105676 597276
rect 105740 597274 105746 597276
rect 106089 597274 106155 597277
rect 105740 597272 106155 597274
rect 105740 597216 106094 597272
rect 106150 597216 106155 597272
rect 105740 597214 106155 597216
rect 105740 597212 105746 597214
rect 106089 597211 106155 597214
rect 230606 597212 230612 597276
rect 230676 597274 230682 597276
rect 231761 597274 231827 597277
rect 230676 597272 231827 597274
rect 230676 597216 231766 597272
rect 231822 597216 231827 597272
rect 230676 597214 231827 597216
rect 230676 597212 230682 597214
rect 231761 597211 231827 597214
rect 422569 597274 422635 597277
rect 422886 597274 422892 597276
rect 422569 597272 422892 597274
rect 422569 597216 422574 597272
rect 422630 597216 422892 597272
rect 422569 597214 422892 597216
rect 422569 597211 422635 597214
rect 422886 597212 422892 597214
rect 422956 597212 422962 597276
rect 426433 597274 426499 597277
rect 427670 597274 427676 597276
rect 426433 597272 427676 597274
rect 426433 597216 426438 597272
rect 426494 597216 427676 597272
rect 426433 597214 427676 597216
rect 426433 597211 426499 597214
rect 427670 597212 427676 597214
rect 427740 597212 427746 597276
rect 427813 597274 427879 597277
rect 428958 597274 428964 597276
rect 427813 597272 428964 597274
rect 427813 597216 427818 597272
rect 427874 597216 428964 597272
rect 427813 597214 428964 597216
rect 427813 597211 427879 597214
rect 428958 597212 428964 597214
rect 429028 597212 429034 597276
rect 430573 597274 430639 597277
rect 430982 597274 430988 597276
rect 430573 597272 430988 597274
rect 430573 597216 430578 597272
rect 430634 597216 430988 597272
rect 430573 597214 430988 597216
rect 430573 597211 430639 597214
rect 430982 597212 430988 597214
rect 431052 597212 431058 597276
rect 99966 597076 99972 597140
rect 100036 597138 100042 597140
rect 100661 597138 100727 597141
rect 104801 597140 104867 597141
rect 100036 597136 100727 597138
rect 100036 597080 100666 597136
rect 100722 597080 100727 597136
rect 100036 597078 100727 597080
rect 100036 597076 100042 597078
rect 100661 597075 100727 597078
rect 104750 597076 104756 597140
rect 104820 597138 104867 597140
rect 204345 597138 204411 597141
rect 205398 597138 205404 597140
rect 104820 597136 104912 597138
rect 104862 597080 104912 597136
rect 104820 597078 104912 597080
rect 204345 597136 205404 597138
rect 204345 597080 204350 597136
rect 204406 597080 205404 597136
rect 204345 597078 205404 597080
rect 104820 597076 104867 597078
rect 104801 597075 104867 597076
rect 204345 597075 204411 597078
rect 205398 597076 205404 597078
rect 205468 597076 205474 597140
rect 349153 597138 349219 597141
rect 350390 597138 350396 597140
rect 349153 597136 350396 597138
rect 349153 597080 349158 597136
rect 349214 597080 350396 597136
rect 349153 597078 350396 597080
rect 349153 597075 349219 597078
rect 350390 597076 350396 597078
rect 350460 597076 350466 597140
rect 429193 597138 429259 597141
rect 429878 597138 429884 597140
rect 429193 597136 429884 597138
rect 429193 597080 429198 597136
rect 429254 597080 429884 597136
rect 429193 597078 429884 597080
rect 429193 597075 429259 597078
rect 429878 597076 429884 597078
rect 429948 597076 429954 597140
rect 94037 597002 94103 597005
rect 94262 597002 94268 597004
rect 94037 597000 94268 597002
rect 94037 596944 94042 597000
rect 94098 596944 94268 597000
rect 94037 596942 94268 596944
rect 94037 596939 94103 596942
rect 94262 596940 94268 596942
rect 94332 596940 94338 597004
rect 97758 596940 97764 597004
rect 97828 597002 97834 597004
rect 97901 597002 97967 597005
rect 97828 597000 97967 597002
rect 97828 596944 97906 597000
rect 97962 596944 97967 597000
rect 97828 596942 97967 596944
rect 97828 596940 97834 596942
rect 97901 596939 97967 596942
rect 130510 596940 130516 597004
rect 130580 597002 130586 597004
rect 131021 597002 131087 597005
rect 130580 597000 131087 597002
rect 130580 596944 131026 597000
rect 131082 596944 131087 597000
rect 130580 596942 131087 596944
rect 130580 596940 130586 596942
rect 131021 596939 131087 596942
rect 314653 597002 314719 597005
rect 315246 597002 315252 597004
rect 314653 597000 315252 597002
rect 314653 596944 314658 597000
rect 314714 596944 315252 597000
rect 314653 596942 315252 596944
rect 314653 596939 314719 596942
rect 315246 596940 315252 596942
rect 315316 596940 315322 597004
rect 339493 597002 339559 597005
rect 340454 597002 340460 597004
rect 339493 597000 340460 597002
rect 339493 596944 339498 597000
rect 339554 596944 340460 597000
rect 339493 596942 340460 596944
rect 339493 596939 339559 596942
rect 340454 596940 340460 596942
rect 340524 596940 340530 597004
rect 423673 597002 423739 597005
rect 424174 597002 424180 597004
rect 423673 597000 424180 597002
rect 423673 596944 423678 597000
rect 423734 596944 424180 597000
rect 423673 596942 424180 596944
rect 423673 596939 423739 596942
rect 424174 596940 424180 596942
rect 424244 596940 424250 597004
rect 431718 596940 431724 597004
rect 431788 597002 431794 597004
rect 431953 597002 432019 597005
rect 433333 597004 433399 597005
rect 434713 597004 434779 597005
rect 433333 597002 433380 597004
rect 431788 597000 432019 597002
rect 431788 596944 431958 597000
rect 432014 596944 432019 597000
rect 431788 596942 432019 596944
rect 433288 597000 433380 597002
rect 433288 596944 433338 597000
rect 433288 596942 433380 596944
rect 431788 596940 431794 596942
rect 431953 596939 432019 596942
rect 433333 596940 433380 596942
rect 433444 596940 433450 597004
rect 434662 596940 434668 597004
rect 434732 597002 434779 597004
rect 434732 597000 434824 597002
rect 434774 596944 434824 597000
rect 434732 596942 434824 596944
rect 434732 596940 434779 596942
rect 433333 596939 433399 596940
rect 434713 596939 434779 596940
rect 110454 596804 110460 596868
rect 110524 596866 110530 596868
rect 173249 596866 173315 596869
rect 110524 596864 173315 596866
rect 110524 596808 173254 596864
rect 173310 596808 173315 596864
rect 110524 596806 173315 596808
rect 110524 596804 110530 596806
rect 173249 596803 173315 596806
rect 240542 596804 240548 596868
rect 240612 596866 240618 596868
rect 241421 596866 241487 596869
rect 240612 596864 241487 596866
rect 240612 596808 241426 596864
rect 241482 596808 241487 596864
rect 240612 596806 241487 596808
rect 240612 596804 240618 596806
rect 241421 596803 241487 596806
rect 313273 596866 313339 596869
rect 314326 596866 314332 596868
rect 313273 596864 314332 596866
rect 313273 596808 313278 596864
rect 313334 596808 314332 596864
rect 313273 596806 314332 596808
rect 313273 596803 313339 596806
rect 314326 596804 314332 596806
rect 314396 596804 314402 596868
rect 409413 596866 409479 596869
rect 465390 596866 465396 596868
rect 409413 596864 465396 596866
rect 409413 596808 409418 596864
rect 409474 596808 465396 596864
rect 409413 596806 465396 596808
rect 409413 596803 409479 596806
rect 465390 596804 465396 596806
rect 465460 596804 465466 596868
rect 125542 596668 125548 596732
rect 125612 596730 125618 596732
rect 126881 596730 126947 596733
rect 125612 596728 126947 596730
rect 125612 596672 126886 596728
rect 126942 596672 126947 596728
rect 125612 596670 126947 596672
rect 125612 596668 125618 596670
rect 126881 596667 126947 596670
rect 434713 596730 434779 596733
rect 435214 596730 435220 596732
rect 434713 596728 435220 596730
rect 434713 596672 434718 596728
rect 434774 596672 435220 596728
rect 434713 596670 435220 596672
rect 434713 596667 434779 596670
rect 435214 596668 435220 596670
rect 435284 596668 435290 596732
rect 444373 596730 444439 596733
rect 445518 596730 445524 596732
rect 444373 596728 445524 596730
rect 444373 596672 444378 596728
rect 444434 596672 445524 596728
rect 444373 596670 445524 596672
rect 444373 596667 444439 596670
rect 445518 596668 445524 596670
rect 445588 596668 445594 596732
rect 135478 596532 135484 596596
rect 135548 596594 135554 596596
rect 136541 596594 136607 596597
rect 140681 596596 140747 596597
rect 135548 596592 136607 596594
rect 135548 596536 136546 596592
rect 136602 596536 136607 596592
rect 135548 596534 136607 596536
rect 135548 596532 135554 596534
rect 136541 596531 136607 596534
rect 140630 596532 140636 596596
rect 140700 596594 140747 596596
rect 311893 596594 311959 596597
rect 312854 596594 312860 596596
rect 140700 596592 140792 596594
rect 140742 596536 140792 596592
rect 140700 596534 140792 596536
rect 311893 596592 312860 596594
rect 311893 596536 311898 596592
rect 311954 596536 312860 596592
rect 311893 596534 312860 596536
rect 140700 596532 140747 596534
rect 140681 596531 140747 596532
rect 311893 596531 311959 596534
rect 312854 596532 312860 596534
rect 312924 596532 312930 596596
rect 202873 596460 202939 596461
rect 202822 596396 202828 596460
rect 202892 596458 202939 596460
rect 425053 596458 425119 596461
rect 425278 596458 425284 596460
rect 202892 596456 202984 596458
rect 202934 596400 202984 596456
rect 202892 596398 202984 596400
rect 425053 596456 425284 596458
rect 425053 596400 425058 596456
rect 425114 596400 425284 596456
rect 425053 596398 425284 596400
rect 202892 596396 202939 596398
rect 202873 596395 202939 596396
rect 425053 596395 425119 596398
rect 425278 596396 425284 596398
rect 425348 596396 425354 596460
rect 95233 596322 95299 596325
rect 95366 596322 95372 596324
rect 95233 596320 95372 596322
rect 95233 596264 95238 596320
rect 95294 596264 95372 596320
rect 95233 596262 95372 596264
rect 95233 596259 95299 596262
rect 95366 596260 95372 596262
rect 95436 596260 95442 596324
rect 115606 596260 115612 596324
rect 115676 596322 115682 596324
rect 115841 596322 115907 596325
rect 115676 596320 115907 596322
rect 115676 596264 115846 596320
rect 115902 596264 115907 596320
rect 115676 596262 115907 596264
rect 115676 596260 115682 596262
rect 115841 596259 115907 596262
rect 120574 596260 120580 596324
rect 120644 596322 120650 596324
rect 121361 596322 121427 596325
rect 204253 596324 204319 596325
rect 204253 596322 204300 596324
rect 120644 596320 121427 596322
rect 120644 596264 121366 596320
rect 121422 596264 121427 596320
rect 120644 596262 121427 596264
rect 204208 596320 204300 596322
rect 204208 596264 204258 596320
rect 204208 596262 204300 596264
rect 120644 596260 120650 596262
rect 121361 596259 121427 596262
rect 204253 596260 204300 596262
rect 204364 596260 204370 596324
rect 219198 596260 219204 596324
rect 219268 596322 219274 596324
rect 219433 596322 219499 596325
rect 219268 596320 219499 596322
rect 219268 596264 219438 596320
rect 219494 596264 219499 596320
rect 219268 596262 219499 596264
rect 219268 596260 219274 596262
rect 204253 596259 204319 596260
rect 219433 596259 219499 596262
rect 335118 596260 335124 596324
rect 335188 596322 335194 596324
rect 335353 596322 335419 596325
rect 335188 596320 335419 596322
rect 335188 596264 335358 596320
rect 335414 596264 335419 596320
rect 335188 596262 335419 596264
rect 335188 596260 335194 596262
rect 335353 596259 335419 596262
rect 354438 596260 354444 596324
rect 354508 596322 354514 596324
rect 354673 596322 354739 596325
rect 455413 596324 455479 596325
rect 455413 596322 455460 596324
rect 354508 596320 354739 596322
rect 354508 596264 354678 596320
rect 354734 596264 354739 596320
rect 354508 596262 354739 596264
rect 455368 596320 455460 596322
rect 455368 596264 455418 596320
rect 455368 596262 455460 596264
rect 354508 596260 354514 596262
rect 354673 596259 354739 596262
rect 455413 596260 455460 596262
rect 455524 596260 455530 596324
rect 470358 596260 470364 596324
rect 470428 596322 470434 596324
rect 470593 596322 470659 596325
rect 470428 596320 470659 596322
rect 470428 596264 470598 596320
rect 470654 596264 470659 596320
rect 470428 596262 470659 596264
rect 470428 596260 470434 596262
rect 455413 596259 455479 596260
rect 470593 596259 470659 596262
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 282126 589868 282132 589932
rect 282196 589930 282202 589932
rect 470593 589930 470659 589933
rect 282196 589928 470659 589930
rect 282196 589872 470598 589928
rect 470654 589872 470659 589928
rect 282196 589870 470659 589872
rect 282196 589868 282202 589870
rect 470593 589867 470659 589870
rect -960 580002 480 580092
rect 3969 580002 4035 580005
rect -960 580000 4035 580002
rect -960 579944 3974 580000
rect 4030 579944 4035 580000
rect -960 579942 4035 579944
rect -960 579852 480 579942
rect 3969 579939 4035 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 187325 527098 187391 527101
rect 298001 527098 298067 527101
rect 187325 527096 189458 527098
rect 187325 527040 187330 527096
rect 187386 527060 189458 527096
rect 298001 527096 299490 527098
rect 187386 527040 190072 527060
rect 187325 527038 190072 527040
rect 187325 527035 187391 527038
rect 78489 526690 78555 526693
rect 80002 526690 80062 527030
rect 189398 527000 190072 527038
rect 298001 527040 298006 527096
rect 298062 527060 299490 527096
rect 298062 527040 300012 527060
rect 298001 527038 300012 527040
rect 298001 527035 298067 527038
rect 299430 527000 300012 527038
rect 78489 526688 80062 526690
rect 78489 526632 78494 526688
rect 78550 526632 80062 526688
rect 78489 526630 80062 526632
rect 78489 526627 78555 526630
rect 407798 526628 407804 526692
rect 407868 526690 407874 526692
rect 410002 526690 410062 527030
rect 407868 526630 410062 526690
rect 407868 526628 407874 526630
rect 78305 526554 78371 526557
rect 407665 526554 407731 526557
rect 78305 526552 80062 526554
rect 78305 526496 78310 526552
rect 78366 526496 80062 526552
rect 78305 526494 80062 526496
rect 78305 526491 78371 526494
rect 80002 525942 80062 526494
rect 407665 526552 410062 526554
rect 407665 526496 407670 526552
rect 407726 526496 410062 526552
rect 407665 526494 410062 526496
rect 407665 526491 407731 526494
rect 186773 526010 186839 526013
rect 188429 526010 188495 526013
rect 297173 526010 297239 526013
rect 186773 526008 189458 526010
rect 186773 525952 186778 526008
rect 186834 525952 188434 526008
rect 188490 525972 189458 526008
rect 297173 526008 299490 526010
rect 188490 525952 190072 525972
rect 186773 525950 190072 525952
rect 186773 525947 186839 525950
rect 188429 525947 188495 525950
rect 189398 525912 190072 525950
rect 297173 525952 297178 526008
rect 297234 525972 299490 526008
rect 297234 525952 300012 525972
rect 297173 525950 300012 525952
rect 297173 525947 297239 525950
rect 299430 525912 300012 525950
rect 410002 525942 410062 526494
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 186865 524378 186931 524381
rect 187509 524378 187575 524381
rect 297357 524378 297423 524381
rect 186865 524376 189458 524378
rect 186865 524320 186870 524376
rect 186926 524320 187514 524376
rect 187570 524340 189458 524376
rect 297357 524376 299490 524378
rect 187570 524320 190072 524340
rect 186865 524318 190072 524320
rect 186865 524315 186931 524318
rect 187509 524315 187575 524318
rect 78305 523698 78371 523701
rect 80002 523698 80062 524310
rect 189398 524280 190072 524318
rect 297357 524320 297362 524376
rect 297418 524340 299490 524376
rect 583520 524364 584960 524454
rect 297418 524320 300012 524340
rect 297357 524318 300012 524320
rect 297357 524315 297423 524318
rect 299430 524280 300012 524318
rect 78305 523696 80062 523698
rect 78305 523640 78310 523696
rect 78366 523640 80062 523696
rect 78305 523638 80062 523640
rect 78305 523635 78371 523638
rect 407614 523636 407620 523700
rect 407684 523698 407690 523700
rect 410002 523698 410062 524310
rect 407684 523638 410062 523698
rect 407684 523636 407690 523638
rect 77753 523562 77819 523565
rect 407757 523562 407823 523565
rect 77753 523560 80062 523562
rect 77753 523504 77758 523560
rect 77814 523504 80062 523560
rect 77753 523502 80062 523504
rect 77753 523499 77819 523502
rect 80002 523222 80062 523502
rect 407757 523560 410062 523562
rect 407757 523504 407762 523560
rect 407818 523504 410062 523560
rect 407757 523502 410062 523504
rect 407757 523499 407823 523502
rect 187417 523290 187483 523293
rect 297633 523290 297699 523293
rect 187417 523288 189458 523290
rect 187417 523232 187422 523288
rect 187478 523252 189458 523288
rect 297633 523288 299490 523290
rect 187478 523232 190072 523252
rect 187417 523230 190072 523232
rect 187417 523227 187483 523230
rect 189398 523192 190072 523230
rect 297633 523232 297638 523288
rect 297694 523252 299490 523288
rect 297694 523232 300012 523252
rect 297633 523230 300012 523232
rect 297633 523227 297699 523230
rect 299430 523192 300012 523230
rect 410002 523222 410062 523502
rect 187233 521658 187299 521661
rect 297265 521658 297331 521661
rect 297725 521658 297791 521661
rect 187233 521656 189458 521658
rect 187233 521600 187238 521656
rect 187294 521620 189458 521656
rect 297265 521656 297791 521658
rect 187294 521600 190072 521620
rect 187233 521598 190072 521600
rect 187233 521595 187299 521598
rect 78121 520978 78187 520981
rect 80002 520978 80062 521590
rect 189398 521560 190072 521598
rect 297265 521600 297270 521656
rect 297326 521600 297730 521656
rect 297786 521600 297791 521656
rect 407481 521658 407547 521661
rect 408217 521658 408283 521661
rect 407481 521656 408283 521658
rect 297265 521598 297791 521600
rect 297265 521595 297331 521598
rect 297725 521595 297791 521598
rect 299798 521560 300012 521620
rect 407481 521600 407486 521656
rect 407542 521600 408222 521656
rect 408278 521600 408283 521656
rect 407481 521598 408283 521600
rect 407481 521595 407547 521598
rect 408217 521595 408283 521598
rect 296805 521522 296871 521525
rect 297449 521522 297515 521525
rect 299798 521522 299858 521560
rect 296805 521520 299858 521522
rect 296805 521464 296810 521520
rect 296866 521464 297454 521520
rect 297510 521464 299858 521520
rect 296805 521462 299858 521464
rect 296805 521459 296871 521462
rect 297449 521459 297515 521462
rect 78121 520976 80062 520978
rect 78121 520920 78126 520976
rect 78182 520920 80062 520976
rect 78121 520918 80062 520920
rect 407665 520978 407731 520981
rect 410002 520978 410062 521590
rect 407665 520976 410062 520978
rect 407665 520920 407670 520976
rect 407726 520920 410062 520976
rect 407665 520918 410062 520920
rect 78121 520915 78187 520918
rect 407665 520915 407731 520918
rect 77845 520298 77911 520301
rect 186681 520298 186747 520301
rect 297265 520298 297331 520301
rect 407481 520298 407547 520301
rect 77845 520296 80062 520298
rect 77845 520240 77850 520296
rect 77906 520240 80062 520296
rect 77845 520238 80062 520240
rect 77845 520235 77911 520238
rect 80002 520230 80062 520238
rect 186681 520296 190010 520298
rect 186681 520240 186686 520296
rect 186742 520260 190010 520296
rect 297265 520296 299858 520298
rect 186742 520240 190072 520260
rect 186681 520238 190072 520240
rect 186681 520235 186747 520238
rect 189950 520200 190072 520238
rect 297265 520240 297270 520296
rect 297326 520260 299858 520296
rect 407481 520296 410062 520298
rect 297326 520240 300012 520260
rect 297265 520238 300012 520240
rect 297265 520235 297331 520238
rect 299798 520200 300012 520238
rect 407481 520240 407486 520296
rect 407542 520240 410062 520296
rect 407481 520238 410062 520240
rect 407481 520235 407547 520238
rect 410002 520230 410062 520238
rect 187141 518666 187207 518669
rect 297541 518666 297607 518669
rect 187141 518664 189458 518666
rect 187141 518608 187146 518664
rect 187202 518628 189458 518664
rect 297541 518664 299490 518666
rect 187202 518608 190072 518628
rect 187141 518606 190072 518608
rect 187141 518603 187207 518606
rect 78581 517986 78647 517989
rect 80002 517986 80062 518598
rect 189398 518568 190072 518606
rect 297541 518608 297546 518664
rect 297602 518628 299490 518664
rect 297602 518608 300012 518628
rect 297541 518606 300012 518608
rect 297541 518603 297607 518606
rect 299430 518568 300012 518606
rect 78581 517984 80062 517986
rect 78581 517928 78586 517984
rect 78642 517928 80062 517984
rect 78581 517926 80062 517928
rect 407389 517986 407455 517989
rect 410002 517986 410062 518598
rect 407389 517984 410062 517986
rect 407389 517928 407394 517984
rect 407450 517928 410062 517984
rect 407389 517926 410062 517928
rect 78581 517923 78647 517926
rect 407389 517923 407455 517926
rect 186773 517578 186839 517581
rect 187141 517578 187207 517581
rect 186773 517576 187207 517578
rect 186773 517520 186778 517576
rect 186834 517520 187146 517576
rect 187202 517520 187207 517576
rect 186773 517518 187207 517520
rect 186773 517515 186839 517518
rect 187141 517515 187207 517518
rect 297541 517578 297607 517581
rect 298001 517578 298067 517581
rect 297541 517576 298067 517578
rect 297541 517520 297546 517576
rect 297602 517520 298006 517576
rect 298062 517520 298067 517576
rect 297541 517518 298067 517520
rect 297541 517515 297607 517518
rect 298001 517515 298067 517518
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 296989 500850 297055 500853
rect 297909 500850 297975 500853
rect 296989 500848 297975 500850
rect 296989 500792 296994 500848
rect 297050 500792 297914 500848
rect 297970 500792 297975 500848
rect 296989 500790 297975 500792
rect 296989 500787 297055 500790
rect 297909 500787 297975 500790
rect 187049 500306 187115 500309
rect 297909 500306 297975 500309
rect 408309 500306 408375 500309
rect 187049 500304 189458 500306
rect 187049 500248 187054 500304
rect 187110 500268 189458 500304
rect 297909 500304 299490 500306
rect 187110 500248 190072 500268
rect 187049 500246 190072 500248
rect 187049 500243 187115 500246
rect 78029 499898 78095 499901
rect 80002 499898 80062 500238
rect 189398 500208 190072 500246
rect 297909 500248 297914 500304
rect 297970 500268 299490 500304
rect 408309 500304 410062 500306
rect 297970 500248 300012 500268
rect 297909 500246 300012 500248
rect 297909 500243 297975 500246
rect 299430 500208 300012 500246
rect 408309 500248 408314 500304
rect 408370 500248 410062 500304
rect 408309 500246 410062 500248
rect 408309 500243 408375 500246
rect 410002 500238 410062 500246
rect 78029 499896 80062 499898
rect 78029 499840 78034 499896
rect 78090 499840 80062 499896
rect 78029 499838 80062 499840
rect 78029 499835 78095 499838
rect 77937 498674 78003 498677
rect 187601 498674 187667 498677
rect 189073 498674 189139 498677
rect 297081 498674 297147 498677
rect 408401 498674 408467 498677
rect 77937 498672 80062 498674
rect 77937 498616 77942 498672
rect 77998 498616 80062 498672
rect 77937 498614 80062 498616
rect 77937 498611 78003 498614
rect 80002 498606 80062 498614
rect 187601 498672 189458 498674
rect 187601 498616 187606 498672
rect 187662 498616 189078 498672
rect 189134 498636 189458 498672
rect 297081 498672 299490 498674
rect 189134 498616 190072 498636
rect 187601 498614 190072 498616
rect 187601 498611 187667 498614
rect 189073 498611 189139 498614
rect 189398 498576 190072 498614
rect 297081 498616 297086 498672
rect 297142 498636 299490 498672
rect 408401 498672 410062 498674
rect 297142 498616 300012 498636
rect 297081 498614 300012 498616
rect 297081 498611 297147 498614
rect 299430 498576 300012 498614
rect 408401 498616 408406 498672
rect 408462 498616 410062 498672
rect 408401 498614 410062 498616
rect 408401 498611 408467 498614
rect 410002 498606 410062 498614
rect 78397 498402 78463 498405
rect 186957 498402 187023 498405
rect 407849 498402 407915 498405
rect 78397 498400 79426 498402
rect 78397 498344 78402 498400
rect 78458 498364 79426 498400
rect 186957 498400 189458 498402
rect 78458 498344 80032 498364
rect 78397 498342 80032 498344
rect 78397 498339 78463 498342
rect 79366 498304 80032 498342
rect 186957 498344 186962 498400
rect 187018 498364 189458 498400
rect 407849 498400 409522 498402
rect 187018 498344 190072 498364
rect 186957 498342 190072 498344
rect 186957 498339 187023 498342
rect 189398 498304 190072 498342
rect 299430 498304 300012 498364
rect 407849 498344 407854 498400
rect 407910 498364 409522 498400
rect 407910 498344 410032 498364
rect 407849 498342 410032 498344
rect 407849 498339 407915 498342
rect 409462 498304 410032 498342
rect 296897 498266 296963 498269
rect 297817 498266 297883 498269
rect 299430 498266 299490 498304
rect 296897 498264 299490 498266
rect 296897 498208 296902 498264
rect 296958 498208 297822 498264
rect 297878 498208 299490 498264
rect 296897 498206 299490 498208
rect 408217 498266 408283 498269
rect 408401 498266 408467 498269
rect 408217 498264 408467 498266
rect 408217 498208 408222 498264
rect 408278 498208 408406 498264
rect 408462 498208 408467 498264
rect 408217 498206 408467 498208
rect 296897 498203 296963 498206
rect 297817 498203 297883 498206
rect 408217 498203 408283 498206
rect 408401 498203 408467 498206
rect 583520 497844 584960 498084
rect 297357 489834 297423 489837
rect 407614 489834 407620 489836
rect 297357 489832 407620 489834
rect 297357 489776 297362 489832
rect 297418 489776 407620 489832
rect 297357 489774 407620 489776
rect 297357 489771 297423 489774
rect 407614 489772 407620 489774
rect 407684 489772 407690 489836
rect -960 488596 480 488836
rect 92933 488476 92999 488477
rect 94221 488476 94287 488477
rect 95325 488476 95391 488477
rect 97809 488476 97875 488477
rect 98913 488476 98979 488477
rect 100017 488476 100083 488477
rect 101121 488476 101187 488477
rect 102409 488476 102475 488477
rect 104801 488476 104867 488477
rect 105721 488476 105787 488477
rect 92933 488472 92980 488476
rect 93044 488474 93050 488476
rect 92933 488416 92938 488472
rect 92933 488412 92980 488416
rect 93044 488414 93090 488474
rect 94221 488472 94268 488476
rect 94332 488474 94338 488476
rect 94221 488416 94226 488472
rect 93044 488412 93050 488414
rect 94221 488412 94268 488416
rect 94332 488414 94378 488474
rect 95325 488472 95372 488476
rect 95436 488474 95442 488476
rect 97758 488474 97764 488476
rect 95325 488416 95330 488472
rect 94332 488412 94338 488414
rect 95325 488412 95372 488416
rect 95436 488414 95482 488474
rect 97718 488414 97764 488474
rect 97828 488472 97875 488476
rect 98862 488474 98868 488476
rect 97870 488416 97875 488472
rect 95436 488412 95442 488414
rect 97758 488412 97764 488414
rect 97828 488412 97875 488416
rect 98822 488414 98868 488474
rect 98932 488472 98979 488476
rect 99966 488474 99972 488476
rect 98974 488416 98979 488472
rect 98862 488412 98868 488414
rect 98932 488412 98979 488416
rect 99926 488414 99972 488474
rect 100036 488472 100083 488476
rect 101070 488474 101076 488476
rect 100078 488416 100083 488472
rect 99966 488412 99972 488414
rect 100036 488412 100083 488416
rect 101030 488414 101076 488474
rect 101140 488472 101187 488476
rect 102358 488474 102364 488476
rect 101182 488416 101187 488472
rect 101070 488412 101076 488414
rect 101140 488412 101187 488416
rect 102318 488414 102364 488474
rect 102428 488472 102475 488476
rect 104750 488474 104756 488476
rect 102470 488416 102475 488472
rect 102358 488412 102364 488414
rect 102428 488412 102475 488416
rect 104710 488414 104756 488474
rect 104820 488472 104867 488476
rect 105670 488474 105676 488476
rect 104862 488416 104867 488472
rect 104750 488412 104756 488414
rect 104820 488412 104867 488416
rect 105630 488414 105676 488474
rect 105740 488472 105787 488476
rect 105782 488416 105787 488472
rect 105670 488412 105676 488414
rect 105740 488412 105787 488416
rect 204294 488412 204300 488476
rect 204364 488474 204370 488476
rect 204437 488474 204503 488477
rect 214833 488476 214899 488477
rect 214782 488474 214788 488476
rect 204364 488472 204503 488474
rect 204364 488416 204442 488472
rect 204498 488416 204503 488472
rect 204364 488414 204503 488416
rect 214742 488414 214788 488474
rect 214852 488472 214899 488476
rect 214894 488416 214899 488472
rect 204364 488412 204370 488414
rect 92933 488411 92999 488412
rect 94221 488411 94287 488412
rect 95325 488411 95391 488412
rect 97809 488411 97875 488412
rect 98913 488411 98979 488412
rect 100017 488411 100083 488412
rect 101121 488411 101187 488412
rect 102409 488411 102475 488412
rect 104801 488411 104867 488412
rect 105721 488411 105787 488412
rect 204437 488411 204503 488414
rect 214782 488412 214788 488414
rect 214852 488412 214899 488416
rect 214833 488411 214899 488412
rect 314285 488476 314351 488477
rect 315389 488476 315455 488477
rect 314285 488472 314332 488476
rect 314396 488474 314402 488476
rect 314285 488416 314290 488472
rect 314285 488412 314332 488416
rect 314396 488414 314442 488474
rect 315389 488472 315436 488476
rect 315500 488474 315506 488476
rect 322933 488474 322999 488477
rect 323342 488474 323348 488476
rect 315389 488416 315394 488472
rect 314396 488412 314402 488414
rect 315389 488412 315436 488416
rect 315500 488414 315546 488474
rect 322933 488472 323348 488474
rect 322933 488416 322938 488472
rect 322994 488416 323348 488472
rect 322933 488414 323348 488416
rect 315500 488412 315506 488414
rect 314285 488411 314351 488412
rect 315389 488411 315455 488412
rect 322933 488411 322999 488414
rect 323342 488412 323348 488414
rect 323412 488412 323418 488476
rect 422569 488474 422635 488477
rect 422886 488474 422892 488476
rect 422569 488472 422892 488474
rect 422569 488416 422574 488472
rect 422630 488416 422892 488472
rect 422569 488414 422892 488416
rect 422569 488411 422635 488414
rect 422886 488412 422892 488414
rect 422956 488412 422962 488476
rect 423673 488474 423739 488477
rect 424174 488474 424180 488476
rect 423673 488472 424180 488474
rect 423673 488416 423678 488472
rect 423734 488416 424180 488472
rect 423673 488414 424180 488416
rect 423673 488411 423739 488414
rect 424174 488412 424180 488414
rect 424244 488412 424250 488476
rect 425053 488474 425119 488477
rect 425278 488474 425284 488476
rect 425053 488472 425284 488474
rect 425053 488416 425058 488472
rect 425114 488416 425284 488472
rect 425053 488414 425284 488416
rect 425053 488411 425119 488414
rect 425278 488412 425284 488414
rect 425348 488412 425354 488476
rect 211153 488340 211219 488341
rect 211102 488338 211108 488340
rect 211062 488278 211108 488338
rect 211172 488336 211219 488340
rect 211214 488280 211219 488336
rect 211102 488276 211108 488278
rect 211172 488276 211219 488280
rect 213494 488276 213500 488340
rect 213564 488338 213570 488340
rect 213729 488338 213795 488341
rect 213564 488336 213795 488338
rect 213564 488280 213734 488336
rect 213790 488280 213795 488336
rect 213564 488278 213795 488280
rect 213564 488276 213570 488278
rect 211153 488275 211219 488276
rect 213729 488275 213795 488278
rect 215385 488338 215451 488341
rect 215702 488338 215708 488340
rect 215385 488336 215708 488338
rect 215385 488280 215390 488336
rect 215446 488280 215708 488336
rect 215385 488278 215708 488280
rect 215385 488275 215451 488278
rect 215702 488276 215708 488278
rect 215772 488276 215778 488340
rect 296805 488338 296871 488341
rect 407665 488338 407731 488341
rect 296805 488336 407731 488338
rect 296805 488280 296810 488336
rect 296866 488280 407670 488336
rect 407726 488280 407731 488336
rect 296805 488278 407731 488280
rect 296805 488275 296871 488278
rect 407665 488275 407731 488278
rect 465073 488338 465139 488341
rect 465390 488338 465396 488340
rect 465073 488336 465396 488338
rect 465073 488280 465078 488336
rect 465134 488280 465396 488336
rect 465073 488278 465396 488280
rect 465073 488275 465139 488278
rect 465390 488276 465396 488278
rect 465460 488276 465466 488340
rect 105302 488140 105308 488204
rect 105372 488202 105378 488204
rect 105997 488202 106063 488205
rect 105372 488200 106063 488202
rect 105372 488144 106002 488200
rect 106058 488144 106063 488200
rect 105372 488142 106063 488144
rect 105372 488140 105378 488142
rect 105997 488139 106063 488142
rect 110454 488140 110460 488204
rect 110524 488202 110530 488204
rect 111701 488202 111767 488205
rect 110524 488200 111767 488202
rect 110524 488144 111706 488200
rect 111762 488144 111767 488200
rect 110524 488142 111767 488144
rect 110524 488140 110530 488142
rect 111701 488139 111767 488142
rect 202873 488202 202939 488205
rect 203006 488202 203012 488204
rect 202873 488200 203012 488202
rect 202873 488144 202878 488200
rect 202934 488144 203012 488200
rect 202873 488142 203012 488144
rect 202873 488139 202939 488142
rect 203006 488140 203012 488142
rect 203076 488140 203082 488204
rect 298001 488202 298067 488205
rect 407389 488202 407455 488205
rect 298001 488200 407455 488202
rect 298001 488144 298006 488200
rect 298062 488144 407394 488200
rect 407450 488144 407455 488200
rect 298001 488142 407455 488144
rect 298001 488139 298067 488142
rect 407389 488139 407455 488142
rect 429193 488202 429259 488205
rect 429878 488202 429884 488204
rect 429193 488200 429884 488202
rect 429193 488144 429198 488200
rect 429254 488144 429884 488200
rect 429193 488142 429884 488144
rect 429193 488139 429259 488142
rect 429878 488140 429884 488142
rect 429948 488140 429954 488204
rect 103278 488004 103284 488068
rect 103348 488066 103354 488068
rect 103421 488066 103487 488069
rect 103348 488064 103487 488066
rect 103348 488008 103426 488064
rect 103482 488008 103487 488064
rect 103348 488006 103487 488008
rect 103348 488004 103354 488006
rect 103421 488003 103487 488006
rect 293401 488066 293467 488069
rect 407798 488066 407804 488068
rect 293401 488064 407804 488066
rect 293401 488008 293406 488064
rect 293462 488008 407804 488064
rect 293401 488006 407804 488008
rect 293401 488003 293467 488006
rect 407798 488004 407804 488006
rect 407868 488004 407874 488068
rect 312997 487932 313063 487933
rect 312997 487928 313044 487932
rect 313108 487930 313114 487932
rect 312997 487872 313002 487928
rect 312997 487868 313044 487872
rect 313108 487870 313154 487930
rect 313108 487868 313114 487870
rect 312997 487867 313063 487868
rect 427813 487794 427879 487797
rect 428958 487794 428964 487796
rect 427813 487792 428964 487794
rect 427813 487736 427818 487792
rect 427874 487736 428964 487792
rect 427813 487734 428964 487736
rect 427813 487731 427879 487734
rect 428958 487732 428964 487734
rect 429028 487732 429034 487796
rect 426433 487658 426499 487661
rect 427670 487658 427676 487660
rect 426433 487656 427676 487658
rect 426433 487600 426438 487656
rect 426494 487600 427676 487656
rect 426433 487598 427676 487600
rect 426433 487595 426499 487598
rect 427670 487596 427676 487598
rect 427740 487596 427746 487660
rect 434713 487658 434779 487661
rect 435582 487658 435588 487660
rect 434713 487656 435588 487658
rect 434713 487600 434718 487656
rect 434774 487600 435588 487656
rect 434713 487598 435588 487600
rect 434713 487595 434779 487598
rect 435582 487596 435588 487598
rect 435652 487596 435658 487660
rect 211797 487522 211863 487525
rect 212206 487522 212212 487524
rect 211797 487520 212212 487522
rect 211797 487464 211802 487520
rect 211858 487464 212212 487520
rect 211797 487462 212212 487464
rect 211797 487459 211863 487462
rect 212206 487460 212212 487462
rect 212276 487460 212282 487524
rect 320909 487522 320975 487525
rect 321134 487522 321140 487524
rect 320909 487520 321140 487522
rect 320909 487464 320914 487520
rect 320970 487464 321140 487520
rect 320909 487462 321140 487464
rect 320909 487459 320975 487462
rect 321134 487460 321140 487462
rect 321204 487460 321210 487524
rect 324814 487460 324820 487524
rect 324884 487522 324890 487524
rect 324957 487522 325023 487525
rect 324884 487520 325023 487522
rect 324884 487464 324962 487520
rect 325018 487464 325023 487520
rect 324884 487462 325023 487464
rect 324884 487460 324890 487462
rect 324957 487459 325023 487462
rect 430573 487522 430639 487525
rect 430982 487522 430988 487524
rect 430573 487520 430988 487522
rect 430573 487464 430578 487520
rect 430634 487464 430988 487520
rect 430573 487462 430988 487464
rect 430573 487459 430639 487462
rect 430982 487460 430988 487462
rect 431052 487460 431058 487524
rect 432137 487522 432203 487525
rect 433333 487524 433399 487525
rect 432270 487522 432276 487524
rect 432137 487520 432276 487522
rect 432137 487464 432142 487520
rect 432198 487464 432276 487520
rect 432137 487462 432276 487464
rect 432137 487459 432203 487462
rect 432270 487460 432276 487462
rect 432340 487460 432346 487524
rect 433333 487522 433380 487524
rect 433288 487520 433380 487522
rect 433288 487464 433338 487520
rect 433288 487462 433380 487464
rect 433333 487460 433380 487462
rect 433444 487460 433450 487524
rect 434713 487522 434779 487525
rect 434846 487522 434852 487524
rect 434713 487520 434852 487522
rect 434713 487464 434718 487520
rect 434774 487464 434852 487520
rect 434713 487462 434852 487464
rect 433333 487459 433399 487460
rect 434713 487459 434779 487462
rect 434846 487460 434852 487462
rect 434916 487460 434922 487524
rect 209998 487324 210004 487388
rect 210068 487386 210074 487388
rect 210417 487386 210483 487389
rect 210068 487384 210483 487386
rect 210068 487328 210422 487384
rect 210478 487328 210483 487384
rect 210068 487326 210483 487328
rect 210068 487324 210074 487326
rect 210417 487323 210483 487326
rect 318926 487324 318932 487388
rect 318996 487386 319002 487388
rect 319621 487386 319687 487389
rect 318996 487384 319687 487386
rect 318996 487328 319626 487384
rect 319682 487328 319687 487384
rect 318996 487326 319687 487328
rect 318996 487324 319002 487326
rect 319621 487323 319687 487326
rect 115606 487188 115612 487252
rect 115676 487250 115682 487252
rect 115841 487250 115907 487253
rect 115676 487248 115907 487250
rect 115676 487192 115846 487248
rect 115902 487192 115907 487248
rect 115676 487190 115907 487192
rect 115676 487188 115682 487190
rect 115841 487187 115907 487190
rect 120574 487188 120580 487252
rect 120644 487250 120650 487252
rect 121361 487250 121427 487253
rect 120644 487248 121427 487250
rect 120644 487192 121366 487248
rect 121422 487192 121427 487248
rect 120644 487190 121427 487192
rect 120644 487188 120650 487190
rect 121361 487187 121427 487190
rect 125542 487188 125548 487252
rect 125612 487250 125618 487252
rect 126881 487250 126947 487253
rect 125612 487248 126947 487250
rect 125612 487192 126886 487248
rect 126942 487192 126947 487248
rect 125612 487190 126947 487192
rect 125612 487188 125618 487190
rect 126881 487187 126947 487190
rect 130510 487188 130516 487252
rect 130580 487250 130586 487252
rect 131021 487250 131087 487253
rect 130580 487248 131087 487250
rect 130580 487192 131026 487248
rect 131082 487192 131087 487248
rect 130580 487190 131087 487192
rect 130580 487188 130586 487190
rect 131021 487187 131087 487190
rect 135478 487188 135484 487252
rect 135548 487250 135554 487252
rect 136541 487250 136607 487253
rect 140681 487252 140747 487253
rect 140630 487250 140636 487252
rect 135548 487248 136607 487250
rect 135548 487192 136546 487248
rect 136602 487192 136607 487248
rect 135548 487190 136607 487192
rect 140590 487190 140636 487250
rect 140700 487248 140747 487252
rect 140742 487192 140747 487248
rect 135548 487188 135554 487190
rect 136541 487187 136607 487190
rect 140630 487188 140636 487190
rect 140700 487188 140747 487192
rect 203006 487188 203012 487252
rect 203076 487250 203082 487252
rect 203517 487250 203583 487253
rect 203076 487248 203583 487250
rect 203076 487192 203522 487248
rect 203578 487192 203583 487248
rect 203076 487190 203583 487192
rect 203076 487188 203082 487190
rect 140681 487187 140747 487188
rect 203517 487187 203583 487190
rect 204897 487250 204963 487253
rect 207657 487252 207723 487253
rect 205398 487250 205404 487252
rect 204897 487248 205404 487250
rect 204897 487192 204902 487248
rect 204958 487192 205404 487248
rect 204897 487190 205404 487192
rect 204897 487187 204963 487190
rect 205398 487188 205404 487190
rect 205468 487188 205474 487252
rect 207606 487250 207612 487252
rect 207566 487190 207612 487250
rect 207676 487248 207723 487252
rect 207718 487192 207723 487248
rect 207606 487188 207612 487190
rect 207676 487188 207723 487192
rect 208894 487188 208900 487252
rect 208964 487250 208970 487252
rect 209037 487250 209103 487253
rect 208964 487248 209103 487250
rect 208964 487192 209042 487248
rect 209098 487192 209103 487248
rect 208964 487190 209103 487192
rect 208964 487188 208970 487190
rect 207657 487187 207723 487188
rect 209037 487187 209103 487190
rect 215334 487188 215340 487252
rect 215404 487250 215410 487252
rect 216581 487250 216647 487253
rect 215404 487248 216647 487250
rect 215404 487192 216586 487248
rect 216642 487192 216647 487248
rect 215404 487190 216647 487192
rect 215404 487188 215410 487190
rect 216581 487187 216647 487190
rect 220486 487188 220492 487252
rect 220556 487250 220562 487252
rect 220721 487250 220787 487253
rect 220556 487248 220787 487250
rect 220556 487192 220726 487248
rect 220782 487192 220787 487248
rect 220556 487190 220787 487192
rect 220556 487188 220562 487190
rect 220721 487187 220787 487190
rect 225454 487188 225460 487252
rect 225524 487250 225530 487252
rect 226241 487250 226307 487253
rect 225524 487248 226307 487250
rect 225524 487192 226246 487248
rect 226302 487192 226307 487248
rect 225524 487190 226307 487192
rect 225524 487188 225530 487190
rect 226241 487187 226307 487190
rect 230606 487188 230612 487252
rect 230676 487250 230682 487252
rect 231761 487250 231827 487253
rect 230676 487248 231827 487250
rect 230676 487192 231766 487248
rect 231822 487192 231827 487248
rect 230676 487190 231827 487192
rect 230676 487188 230682 487190
rect 231761 487187 231827 487190
rect 235574 487188 235580 487252
rect 235644 487250 235650 487252
rect 235901 487250 235967 487253
rect 235644 487248 235967 487250
rect 235644 487192 235906 487248
rect 235962 487192 235967 487248
rect 235644 487190 235967 487192
rect 235644 487188 235650 487190
rect 235901 487187 235967 487190
rect 240542 487188 240548 487252
rect 240612 487250 240618 487252
rect 241421 487250 241487 487253
rect 240612 487248 241487 487250
rect 240612 487192 241426 487248
rect 241482 487192 241487 487248
rect 240612 487190 241487 487192
rect 240612 487188 240618 487190
rect 241421 487187 241487 487190
rect 244641 487250 244707 487253
rect 245510 487250 245516 487252
rect 244641 487248 245516 487250
rect 244641 487192 244646 487248
rect 244702 487192 245516 487248
rect 244641 487190 245516 487192
rect 244641 487187 244707 487190
rect 245510 487188 245516 487190
rect 245580 487188 245586 487252
rect 249977 487250 250043 487253
rect 250478 487250 250484 487252
rect 249977 487248 250484 487250
rect 249977 487192 249982 487248
rect 250038 487192 250484 487248
rect 249977 487190 250484 487192
rect 249977 487187 250043 487190
rect 250478 487188 250484 487190
rect 250548 487188 250554 487252
rect 317638 487188 317644 487252
rect 317708 487250 317714 487252
rect 318057 487250 318123 487253
rect 317708 487248 318123 487250
rect 317708 487192 318062 487248
rect 318118 487192 318123 487248
rect 317708 487190 318123 487192
rect 317708 487188 317714 487190
rect 318057 487187 318123 487190
rect 319437 487250 319503 487253
rect 320081 487252 320147 487253
rect 320030 487250 320036 487252
rect 319437 487248 320036 487250
rect 320100 487250 320147 487252
rect 322197 487252 322263 487253
rect 320100 487248 320228 487250
rect 319437 487192 319442 487248
rect 319498 487192 320036 487248
rect 320142 487192 320228 487248
rect 319437 487190 320036 487192
rect 319437 487187 319503 487190
rect 320030 487188 320036 487190
rect 320100 487190 320228 487192
rect 322197 487248 322244 487252
rect 322308 487250 322314 487252
rect 324313 487250 324379 487253
rect 325182 487250 325188 487252
rect 322197 487192 322202 487248
rect 320100 487188 320147 487190
rect 320081 487187 320147 487188
rect 322197 487188 322244 487192
rect 322308 487190 322354 487250
rect 324313 487248 325188 487250
rect 324313 487192 324318 487248
rect 324374 487192 325188 487248
rect 324313 487190 325188 487192
rect 322308 487188 322314 487190
rect 322197 487187 322263 487188
rect 324313 487187 324379 487190
rect 325182 487188 325188 487190
rect 325252 487188 325258 487252
rect 325734 487188 325740 487252
rect 325804 487250 325810 487252
rect 326337 487250 326403 487253
rect 325804 487248 326403 487250
rect 325804 487192 326342 487248
rect 326398 487192 326403 487248
rect 325804 487190 326403 487192
rect 325804 487188 325810 487190
rect 326337 487187 326403 487190
rect 329833 487250 329899 487253
rect 330518 487250 330524 487252
rect 329833 487248 330524 487250
rect 329833 487192 329838 487248
rect 329894 487192 330524 487248
rect 329833 487190 330524 487192
rect 329833 487187 329899 487190
rect 330518 487188 330524 487190
rect 330588 487188 330594 487252
rect 335353 487250 335419 487253
rect 335486 487250 335492 487252
rect 335353 487248 335492 487250
rect 335353 487192 335358 487248
rect 335414 487192 335492 487248
rect 335353 487190 335492 487192
rect 335353 487187 335419 487190
rect 335486 487188 335492 487190
rect 335556 487188 335562 487252
rect 339493 487250 339559 487253
rect 340454 487250 340460 487252
rect 339493 487248 340460 487250
rect 339493 487192 339498 487248
rect 339554 487192 340460 487248
rect 339493 487190 340460 487192
rect 339493 487187 339559 487190
rect 340454 487188 340460 487190
rect 340524 487188 340530 487252
rect 345013 487250 345079 487253
rect 345606 487250 345612 487252
rect 345013 487248 345612 487250
rect 345013 487192 345018 487248
rect 345074 487192 345612 487248
rect 345013 487190 345612 487192
rect 345013 487187 345079 487190
rect 345606 487188 345612 487190
rect 345676 487188 345682 487252
rect 349153 487250 349219 487253
rect 350390 487250 350396 487252
rect 349153 487248 350396 487250
rect 349153 487192 349158 487248
rect 349214 487192 350396 487248
rect 349153 487190 350396 487192
rect 349153 487187 349219 487190
rect 350390 487188 350396 487190
rect 350460 487188 350466 487252
rect 354673 487250 354739 487253
rect 355542 487250 355548 487252
rect 354673 487248 355548 487250
rect 354673 487192 354678 487248
rect 354734 487192 355548 487248
rect 354673 487190 355548 487192
rect 354673 487187 354739 487190
rect 355542 487188 355548 487190
rect 355612 487188 355618 487252
rect 360193 487250 360259 487253
rect 360510 487250 360516 487252
rect 360193 487248 360516 487250
rect 360193 487192 360198 487248
rect 360254 487192 360516 487248
rect 360193 487190 360516 487192
rect 360193 487187 360259 487190
rect 360510 487188 360516 487190
rect 360580 487188 360586 487252
rect 434713 487250 434779 487253
rect 435214 487250 435220 487252
rect 434713 487248 435220 487250
rect 434713 487192 434718 487248
rect 434774 487192 435220 487248
rect 434713 487190 435220 487192
rect 434713 487187 434779 487190
rect 435214 487188 435220 487190
rect 435284 487188 435290 487252
rect 440233 487250 440299 487253
rect 440366 487250 440372 487252
rect 440233 487248 440372 487250
rect 440233 487192 440238 487248
rect 440294 487192 440372 487248
rect 440233 487190 440372 487192
rect 440233 487187 440299 487190
rect 440366 487188 440372 487190
rect 440436 487188 440442 487252
rect 444373 487250 444439 487253
rect 445518 487250 445524 487252
rect 444373 487248 445524 487250
rect 444373 487192 444378 487248
rect 444434 487192 445524 487248
rect 444373 487190 445524 487192
rect 444373 487187 444439 487190
rect 445518 487188 445524 487190
rect 445588 487188 445594 487252
rect 449893 487250 449959 487253
rect 450486 487250 450492 487252
rect 449893 487248 450492 487250
rect 449893 487192 449898 487248
rect 449954 487192 450492 487248
rect 449893 487190 450492 487192
rect 449893 487187 449959 487190
rect 450486 487188 450492 487190
rect 450556 487188 450562 487252
rect 454677 487250 454743 487253
rect 455454 487250 455460 487252
rect 454677 487248 455460 487250
rect 454677 487192 454682 487248
rect 454738 487192 455460 487248
rect 454677 487190 455460 487192
rect 454677 487187 454743 487190
rect 455454 487188 455460 487190
rect 455524 487188 455530 487252
rect 459553 487250 459619 487253
rect 460422 487250 460428 487252
rect 459553 487248 460428 487250
rect 459553 487192 459558 487248
rect 459614 487192 460428 487248
rect 459553 487190 460428 487192
rect 459553 487187 459619 487190
rect 460422 487188 460428 487190
rect 460492 487188 460498 487252
rect 470593 487250 470659 487253
rect 470726 487250 470732 487252
rect 470593 487248 470732 487250
rect 470593 487192 470598 487248
rect 470654 487192 470732 487248
rect 470593 487190 470732 487192
rect 470593 487187 470659 487190
rect 470726 487188 470732 487190
rect 470796 487188 470802 487252
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2865 462634 2931 462637
rect -960 462632 2931 462634
rect -960 462576 2870 462632
rect 2926 462576 2931 462632
rect -960 462574 2931 462576
rect -960 462484 480 462574
rect 2865 462571 2931 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 232129 454338 232195 454341
rect 382222 454338 382228 454340
rect 232129 454336 382228 454338
rect 232129 454280 232134 454336
rect 232190 454280 382228 454336
rect 232129 454278 382228 454280
rect 232129 454275 232195 454278
rect 382222 454276 382228 454278
rect 382292 454276 382298 454340
rect 232681 454202 232747 454205
rect 378726 454202 378732 454204
rect 232681 454200 378732 454202
rect 232681 454144 232686 454200
rect 232742 454144 378732 454200
rect 232681 454142 378732 454144
rect 232681 454139 232747 454142
rect 378726 454140 378732 454142
rect 378796 454140 378802 454204
rect 383929 454202 383995 454205
rect 378918 454200 383995 454202
rect 378918 454144 383934 454200
rect 383990 454144 383995 454200
rect 378918 454142 383995 454144
rect 225689 454066 225755 454069
rect 225689 454064 378610 454066
rect 225689 454008 225694 454064
rect 225750 454008 378610 454064
rect 225689 454006 378610 454008
rect 225689 454003 225755 454006
rect 378550 453930 378610 454006
rect 378918 453930 378978 454142
rect 383929 454139 383995 454142
rect 379094 454004 379100 454068
rect 379164 454066 379170 454068
rect 385125 454066 385191 454069
rect 379164 454064 385191 454066
rect 379164 454008 385130 454064
rect 385186 454008 385191 454064
rect 379164 454006 385191 454008
rect 379164 454004 379170 454006
rect 385125 454003 385191 454006
rect 378550 453870 378978 453930
rect 297817 452434 297883 452437
rect 297817 452432 300196 452434
rect 297817 452376 297822 452432
rect 297878 452376 300196 452432
rect 297817 452374 300196 452376
rect 297817 452371 297883 452374
rect 384021 452298 384087 452301
rect 383886 452296 384087 452298
rect 383886 452240 384026 452296
rect 384082 452240 384087 452296
rect 383886 452238 384087 452240
rect 383886 451724 383946 452238
rect 384021 452235 384087 452238
rect 234061 449850 234127 449853
rect 297357 449850 297423 449853
rect 234061 449848 297423 449850
rect 234061 449792 234066 449848
rect 234122 449792 297362 449848
rect 297418 449792 297423 449848
rect 234061 449790 297423 449792
rect 234061 449787 234127 449790
rect 297357 449787 297423 449790
rect 234245 449714 234311 449717
rect 234521 449714 234587 449717
rect 297173 449714 297239 449717
rect 234245 449712 297239 449714
rect -960 449578 480 449668
rect 234245 449656 234250 449712
rect 234306 449656 234526 449712
rect 234582 449656 297178 449712
rect 297234 449656 297239 449712
rect 234245 449654 297239 449656
rect 234245 449651 234311 449654
rect 234521 449651 234587 449654
rect 297173 449651 297239 449654
rect 3233 449578 3299 449581
rect -960 449576 3299 449578
rect -960 449520 3238 449576
rect 3294 449520 3299 449576
rect -960 449518 3299 449520
rect -960 449428 480 449518
rect 3233 449515 3299 449518
rect 255405 449578 255471 449581
rect 256417 449578 256483 449581
rect 291929 449578 291995 449581
rect 255405 449576 291995 449578
rect 255405 449520 255410 449576
rect 255466 449520 256422 449576
rect 256478 449520 291934 449576
rect 291990 449520 291995 449576
rect 255405 449518 291995 449520
rect 255405 449515 255471 449518
rect 256417 449515 256483 449518
rect 291929 449515 291995 449518
rect 224401 448626 224467 448629
rect 299381 448626 299447 448629
rect 224401 448624 299447 448626
rect 224401 448568 224406 448624
rect 224462 448568 299386 448624
rect 299442 448568 299447 448624
rect 224401 448566 299447 448568
rect 224401 448563 224467 448566
rect 299381 448563 299447 448566
rect 298001 448354 298067 448357
rect 298001 448352 300196 448354
rect 298001 448296 298006 448352
rect 298062 448296 300196 448352
rect 298001 448294 300196 448296
rect 298001 448291 298067 448294
rect 384021 448218 384087 448221
rect 383886 448216 384087 448218
rect 383886 448160 384026 448216
rect 384082 448160 384087 448216
rect 383886 448158 384087 448160
rect 383886 447644 383946 448158
rect 384021 448155 384087 448158
rect 3550 446796 3556 446860
rect 3620 446858 3626 446860
rect 229185 446858 229251 446861
rect 3620 446856 229251 446858
rect 3620 446800 229190 446856
rect 229246 446800 229251 446856
rect 3620 446798 229251 446800
rect 3620 446796 3626 446798
rect 229185 446795 229251 446798
rect 229001 446722 229067 446725
rect 264973 446722 265039 446725
rect 229001 446720 265039 446722
rect 229001 446664 229006 446720
rect 229062 446664 264978 446720
rect 265034 446664 265039 446720
rect 229001 446662 265039 446664
rect 229001 446659 229067 446662
rect 264973 446659 265039 446662
rect 202086 446524 202092 446588
rect 202156 446586 202162 446588
rect 227161 446586 227227 446589
rect 202156 446584 227227 446586
rect 202156 446528 227166 446584
rect 227222 446528 227227 446584
rect 202156 446526 227227 446528
rect 202156 446524 202162 446526
rect 227161 446523 227227 446526
rect 230381 446586 230447 446589
rect 256601 446586 256667 446589
rect 230381 446584 256667 446586
rect 230381 446528 230386 446584
rect 230442 446528 256606 446584
rect 256662 446528 256667 446584
rect 230381 446526 256667 446528
rect 230381 446523 230447 446526
rect 256601 446523 256667 446526
rect 3366 446388 3372 446452
rect 3436 446450 3442 446452
rect 229737 446450 229803 446453
rect 3436 446448 229803 446450
rect 3436 446392 229742 446448
rect 229798 446392 229803 446448
rect 3436 446390 229803 446392
rect 3436 446388 3442 446390
rect 229737 446387 229803 446390
rect 255497 446450 255563 446453
rect 282126 446450 282132 446452
rect 255497 446448 282132 446450
rect 255497 446392 255502 446448
rect 255558 446392 282132 446448
rect 255497 446390 282132 446392
rect 255497 446387 255563 446390
rect 282126 446388 282132 446390
rect 282196 446388 282202 446452
rect 298093 446450 298159 446453
rect 298502 446450 298508 446452
rect 298093 446448 298508 446450
rect 298093 446392 298098 446448
rect 298154 446392 298508 446448
rect 298093 446390 298508 446392
rect 298093 446387 298159 446390
rect 298502 446388 298508 446390
rect 298572 446388 298578 446452
rect 213177 446314 213243 446317
rect 299105 446314 299171 446317
rect 213177 446312 299171 446314
rect 213177 446256 213182 446312
rect 213238 446256 299110 446312
rect 299166 446256 299171 446312
rect 213177 446254 299171 446256
rect 213177 446251 213243 446254
rect 299105 446251 299171 446254
rect 212073 446178 212139 446181
rect 298921 446178 298987 446181
rect 212073 446176 298987 446178
rect 212073 446120 212078 446176
rect 212134 446120 298926 446176
rect 298982 446120 298987 446176
rect 212073 446118 298987 446120
rect 212073 446115 212139 446118
rect 298921 446115 298987 446118
rect 210417 446042 210483 446045
rect 298737 446042 298803 446045
rect 210417 446040 298803 446042
rect 210417 445984 210422 446040
rect 210478 445984 298742 446040
rect 298798 445984 298803 446040
rect 210417 445982 298803 445984
rect 210417 445979 210483 445982
rect 298737 445979 298803 445982
rect 226241 445906 226307 445909
rect 264278 445906 264284 445908
rect 226241 445904 264284 445906
rect 226241 445848 226246 445904
rect 226302 445848 264284 445904
rect 226241 445846 264284 445848
rect 226241 445843 226307 445846
rect 264278 445844 264284 445846
rect 264348 445844 264354 445908
rect 256785 445770 256851 445773
rect 262622 445770 262628 445772
rect 256785 445768 262628 445770
rect 256785 445712 256790 445768
rect 256846 445712 262628 445768
rect 256785 445710 262628 445712
rect 256785 445707 256851 445710
rect 262622 445708 262628 445710
rect 262692 445708 262698 445772
rect 210233 445090 210299 445093
rect 231393 445090 231459 445093
rect 262806 445090 262812 445092
rect 210233 445088 215310 445090
rect 210233 445032 210238 445088
rect 210294 445032 215310 445088
rect 210233 445030 215310 445032
rect 210233 445027 210299 445030
rect 209681 444954 209747 444957
rect 215250 444954 215310 445030
rect 231393 445088 262812 445090
rect 231393 445032 231398 445088
rect 231454 445032 262812 445088
rect 231393 445030 262812 445032
rect 231393 445027 231459 445030
rect 262806 445028 262812 445030
rect 262876 445028 262882 445092
rect 265801 444954 265867 444957
rect 209681 444952 214666 444954
rect 209681 444896 209686 444952
rect 209742 444896 214666 444952
rect 209681 444894 214666 444896
rect 215250 444952 265867 444954
rect 215250 444896 265806 444952
rect 265862 444896 265867 444952
rect 215250 444894 265867 444896
rect 209681 444891 209747 444894
rect 214606 444818 214666 444894
rect 265801 444891 265867 444894
rect 265617 444818 265683 444821
rect 214606 444816 265683 444818
rect 214606 444760 265622 444816
rect 265678 444760 265683 444816
rect 214606 444758 265683 444760
rect 265617 444755 265683 444758
rect 210049 444682 210115 444685
rect 283557 444682 283623 444685
rect 210049 444680 283623 444682
rect 210049 444624 210054 444680
rect 210110 444624 283562 444680
rect 283618 444624 283623 444680
rect 583520 444668 584960 444908
rect 210049 444622 283623 444624
rect 210049 444619 210115 444622
rect 283557 444619 283623 444622
rect 210601 444546 210667 444549
rect 296069 444546 296135 444549
rect 210601 444544 296135 444546
rect 210601 444488 210606 444544
rect 210662 444488 296074 444544
rect 296130 444488 296135 444544
rect 210601 444486 296135 444488
rect 210601 444483 210667 444486
rect 296069 444483 296135 444486
rect 209497 444410 209563 444413
rect 295926 444410 295932 444412
rect 209497 444408 295932 444410
rect 209497 444352 209502 444408
rect 209558 444352 295932 444408
rect 209497 444350 295932 444352
rect 209497 444347 209563 444350
rect 295926 444348 295932 444350
rect 295996 444348 296002 444412
rect 211705 444138 211771 444141
rect 211838 444138 211844 444140
rect 211705 444136 211844 444138
rect 211705 444080 211710 444136
rect 211766 444080 211844 444136
rect 211705 444078 211844 444080
rect 211705 444075 211771 444078
rect 211838 444076 211844 444078
rect 211908 444076 211914 444140
rect 212257 444138 212323 444141
rect 212390 444138 212396 444140
rect 212257 444136 212396 444138
rect 212257 444080 212262 444136
rect 212318 444080 212396 444136
rect 212257 444078 212396 444080
rect 212257 444075 212323 444078
rect 212390 444076 212396 444078
rect 212460 444076 212466 444140
rect 212809 444138 212875 444141
rect 212942 444138 212948 444140
rect 212809 444136 212948 444138
rect 212809 444080 212814 444136
rect 212870 444080 212948 444136
rect 212809 444078 212948 444080
rect 212809 444075 212875 444078
rect 212942 444076 212948 444078
rect 213012 444076 213018 444140
rect 250897 444138 250963 444141
rect 251030 444138 251036 444140
rect 250897 444136 251036 444138
rect 250897 444080 250902 444136
rect 250958 444080 251036 444136
rect 250897 444078 251036 444080
rect 250897 444075 250963 444078
rect 251030 444076 251036 444078
rect 251100 444076 251106 444140
rect 256417 444138 256483 444141
rect 256550 444138 256556 444140
rect 256417 444136 256556 444138
rect 256417 444080 256422 444136
rect 256478 444080 256556 444136
rect 256417 444078 256556 444080
rect 256417 444075 256483 444078
rect 256550 444076 256556 444078
rect 256620 444076 256626 444140
rect 209957 444002 210023 444005
rect 220077 444002 220143 444005
rect 209957 444000 220143 444002
rect 209957 443944 209962 444000
rect 210018 443944 220082 444000
rect 220138 443944 220143 444000
rect 209957 443942 220143 443944
rect 209957 443939 210023 443942
rect 220077 443939 220143 443942
rect 211613 443866 211679 443869
rect 298829 443866 298895 443869
rect 211613 443864 298895 443866
rect 211613 443808 211618 443864
rect 211674 443808 298834 443864
rect 298890 443808 298895 443864
rect 211613 443806 298895 443808
rect 211613 443803 211679 443806
rect 298829 443803 298895 443806
rect 211245 443730 211311 443733
rect 265893 443730 265959 443733
rect 211245 443728 265959 443730
rect 211245 443672 211250 443728
rect 211306 443672 265898 443728
rect 265954 443672 265959 443728
rect 211245 443670 265959 443672
rect 211245 443667 211311 443670
rect 265893 443667 265959 443670
rect 209405 443594 209471 443597
rect 264094 443594 264100 443596
rect 209405 443592 264100 443594
rect 209405 443536 209410 443592
rect 209466 443536 264100 443592
rect 209405 443534 264100 443536
rect 209405 443531 209471 443534
rect 264094 443532 264100 443534
rect 264164 443532 264170 443596
rect 298001 443594 298067 443597
rect 298001 443592 300196 443594
rect 298001 443536 298006 443592
rect 298062 443536 300196 443592
rect 298001 443534 300196 443536
rect 298001 443531 298067 443534
rect 211981 443458 212047 443461
rect 212717 443458 212783 443461
rect 215845 443458 215911 443461
rect 216581 443458 216647 443461
rect 211981 443456 212642 443458
rect 211981 443400 211986 443456
rect 212042 443400 212642 443456
rect 211981 443398 212642 443400
rect 211981 443395 212047 443398
rect 212582 443186 212642 443398
rect 212717 443456 215310 443458
rect 212717 443400 212722 443456
rect 212778 443400 215310 443456
rect 212717 443398 215310 443400
rect 212717 443395 212783 443398
rect 215250 443322 215310 443398
rect 215845 443456 216647 443458
rect 215845 443400 215850 443456
rect 215906 443400 216586 443456
rect 216642 443400 216647 443456
rect 215845 443398 216647 443400
rect 215845 443395 215911 443398
rect 216581 443395 216647 443398
rect 220077 443458 220143 443461
rect 265709 443458 265775 443461
rect 220077 443456 265775 443458
rect 220077 443400 220082 443456
rect 220138 443400 265714 443456
rect 265770 443400 265775 443456
rect 220077 443398 265775 443400
rect 220077 443395 220143 443398
rect 265709 443395 265775 443398
rect 299197 443322 299263 443325
rect 215250 443320 299263 443322
rect 215250 443264 299202 443320
rect 299258 443264 299263 443320
rect 215250 443262 299263 443264
rect 299197 443259 299263 443262
rect 299013 443186 299079 443189
rect 212582 443184 299079 443186
rect 212582 443128 299018 443184
rect 299074 443128 299079 443184
rect 212582 443126 299079 443128
rect 299013 443123 299079 443126
rect 385493 442914 385559 442917
rect 383916 442912 385559 442914
rect 383916 442856 385498 442912
rect 385554 442856 385559 442912
rect 383916 442854 385559 442856
rect 385493 442851 385559 442854
rect 251030 442716 251036 442780
rect 251100 442778 251106 442780
rect 292941 442778 293007 442781
rect 251100 442776 293007 442778
rect 251100 442720 292946 442776
rect 293002 442720 293007 442776
rect 251100 442718 293007 442720
rect 251100 442716 251106 442718
rect 292941 442715 293007 442718
rect 256550 442580 256556 442644
rect 256620 442642 256626 442644
rect 299841 442642 299907 442645
rect 256620 442640 299907 442642
rect 256620 442584 299846 442640
rect 299902 442584 299907 442640
rect 256620 442582 299907 442584
rect 256620 442580 256626 442582
rect 299841 442579 299907 442582
rect 212942 442444 212948 442508
rect 213012 442506 213018 442508
rect 296345 442506 296411 442509
rect 213012 442504 296411 442506
rect 213012 442448 296350 442504
rect 296406 442448 296411 442504
rect 213012 442446 296411 442448
rect 213012 442444 213018 442446
rect 296345 442443 296411 442446
rect 211838 442308 211844 442372
rect 211908 442370 211914 442372
rect 295977 442370 296043 442373
rect 211908 442368 296043 442370
rect 211908 442312 295982 442368
rect 296038 442312 296043 442368
rect 211908 442310 296043 442312
rect 211908 442308 211914 442310
rect 295977 442307 296043 442310
rect 212390 442172 212396 442236
rect 212460 442234 212466 442236
rect 296161 442234 296227 442237
rect 212460 442232 296227 442234
rect 212460 442176 296166 442232
rect 296222 442176 296227 442232
rect 212460 442174 296227 442176
rect 212460 442172 212466 442174
rect 296161 442171 296227 442174
rect 298001 439514 298067 439517
rect 298001 439512 300196 439514
rect 298001 439456 298006 439512
rect 298062 439456 300196 439512
rect 298001 439454 300196 439456
rect 298001 439451 298067 439454
rect 383886 438701 383946 438804
rect 383886 438696 383995 438701
rect 383886 438640 383934 438696
rect 383990 438640 383995 438696
rect 383886 438638 383995 438640
rect 383929 438635 383995 438638
rect -960 436508 480 436748
rect 297173 434754 297239 434757
rect 297173 434752 300196 434754
rect 297173 434696 297178 434752
rect 297234 434696 300196 434752
rect 297173 434694 300196 434696
rect 297173 434691 297239 434694
rect 385401 434074 385467 434077
rect 383916 434072 385467 434074
rect 383916 434016 385406 434072
rect 385462 434016 385467 434072
rect 383916 434014 385467 434016
rect 385401 434011 385467 434014
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 298001 430674 298067 430677
rect 298001 430672 300196 430674
rect 298001 430616 298006 430672
rect 298062 430616 300196 430672
rect 298001 430614 300196 430616
rect 298001 430611 298067 430614
rect 385309 429994 385375 429997
rect 383916 429992 385375 429994
rect 383916 429936 385314 429992
rect 385370 429936 385375 429992
rect 383916 429934 385375 429936
rect 385309 429931 385375 429934
rect 298001 425914 298067 425917
rect 298001 425912 300196 425914
rect 298001 425856 298006 425912
rect 298062 425856 300196 425912
rect 298001 425854 300196 425856
rect 298001 425851 298067 425854
rect 383326 425716 383332 425780
rect 383396 425716 383402 425780
rect 383334 425204 383394 425716
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 297541 421834 297607 421837
rect 297541 421832 300196 421834
rect 297541 421776 297546 421832
rect 297602 421776 300196 421832
rect 297541 421774 300196 421776
rect 297541 421771 297607 421774
rect 383929 421698 383995 421701
rect 383886 421696 383995 421698
rect 383886 421640 383934 421696
rect 383990 421640 383995 421696
rect 383886 421635 383995 421640
rect 383886 421124 383946 421635
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 297449 417074 297515 417077
rect 297449 417072 300196 417074
rect 297449 417016 297454 417072
rect 297510 417016 300196 417072
rect 297449 417014 300196 417016
rect 297449 417011 297515 417014
rect 385217 416394 385283 416397
rect 383916 416392 385283 416394
rect 383916 416336 385222 416392
rect 385278 416336 385283 416392
rect 383916 416334 385283 416336
rect 385217 416331 385283 416334
rect 297357 412994 297423 412997
rect 297357 412992 300196 412994
rect 297357 412936 297362 412992
rect 297418 412936 300196 412992
rect 297357 412934 300196 412936
rect 297357 412931 297423 412934
rect 385125 412314 385191 412317
rect 383916 412312 385191 412314
rect 383916 412256 385130 412312
rect 385186 412256 385191 412312
rect 383916 412254 385191 412256
rect 385125 412251 385191 412254
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 298001 408234 298067 408237
rect 298001 408232 300196 408234
rect 298001 408176 298006 408232
rect 298062 408176 300196 408232
rect 298001 408174 300196 408176
rect 298001 408171 298067 408174
rect 385033 407554 385099 407557
rect 383916 407552 385099 407554
rect 383916 407496 385038 407552
rect 385094 407496 385099 407552
rect 383916 407494 385099 407496
rect 385033 407491 385099 407494
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect 298001 404154 298067 404157
rect 298001 404152 300196 404154
rect 298001 404096 298006 404152
rect 298062 404096 300196 404152
rect 298001 404094 300196 404096
rect 298001 404091 298067 404094
rect 385033 403474 385099 403477
rect 383916 403472 385099 403474
rect 383916 403416 385038 403472
rect 385094 403416 385099 403472
rect 383916 403414 385099 403416
rect 385033 403411 385099 403414
rect 293125 401026 293191 401029
rect 332542 401026 332548 401028
rect 293125 401024 332548 401026
rect 293125 400968 293130 401024
rect 293186 400968 332548 401024
rect 293125 400966 332548 400968
rect 293125 400963 293191 400966
rect 332542 400964 332548 400966
rect 332612 400964 332618 401028
rect 292941 400890 293007 400893
rect 292941 400888 374010 400890
rect 292941 400832 292946 400888
rect 293002 400832 374010 400888
rect 292941 400830 374010 400832
rect 292941 400827 293007 400830
rect 313273 400618 313339 400621
rect 332593 400620 332659 400621
rect 234846 400616 313339 400618
rect 234846 400560 313278 400616
rect 313334 400560 313339 400616
rect 234846 400558 313339 400560
rect 234705 399938 234771 399941
rect 234846 399938 234906 400558
rect 313273 400555 313339 400558
rect 332542 400556 332548 400620
rect 332612 400618 332659 400620
rect 373950 400618 374010 400830
rect 382733 400618 382799 400621
rect 332612 400616 332704 400618
rect 332654 400560 332704 400616
rect 332612 400558 332704 400560
rect 373950 400616 382799 400618
rect 373950 400560 382738 400616
rect 382794 400560 382799 400616
rect 373950 400558 382799 400560
rect 332612 400556 332659 400558
rect 332593 400555 332659 400556
rect 382733 400555 382799 400558
rect 383653 400482 383719 400485
rect 240366 400480 383719 400482
rect 240366 400424 383658 400480
rect 383714 400424 383719 400480
rect 240366 400422 383719 400424
rect 234705 399936 234906 399938
rect 234705 399880 234710 399936
rect 234766 399880 234906 399936
rect 234705 399878 234906 399880
rect 240225 399938 240291 399941
rect 240366 399938 240426 400422
rect 383653 400419 383719 400422
rect 455413 400346 455479 400349
rect 245886 400344 455479 400346
rect 245886 400288 455418 400344
rect 455474 400288 455479 400344
rect 245886 400286 455479 400288
rect 240225 399936 240426 399938
rect 240225 399880 240230 399936
rect 240286 399880 240426 399936
rect 240225 399878 240426 399880
rect 245745 399938 245811 399941
rect 245886 399938 245946 400286
rect 455413 400283 455479 400286
rect 245745 399936 245946 399938
rect 245745 399880 245750 399936
rect 245806 399880 245946 399936
rect 245745 399878 245946 399880
rect 234705 399875 234771 399878
rect 240225 399875 240291 399878
rect 245745 399875 245811 399878
rect 253054 399196 253060 399260
rect 253124 399258 253130 399260
rect 253657 399258 253723 399261
rect 253124 399256 253723 399258
rect 253124 399200 253662 399256
rect 253718 399200 253723 399256
rect 253124 399198 253723 399200
rect 253124 399196 253130 399198
rect 253657 399195 253723 399198
rect 219341 399122 219407 399125
rect 219206 399120 219407 399122
rect 219206 399064 219346 399120
rect 219402 399064 219407 399120
rect 219206 399062 219407 399064
rect 207749 398850 207815 398853
rect 214005 398850 214071 398853
rect 217225 398850 217291 398853
rect 207749 398848 214071 398850
rect 207749 398792 207754 398848
rect 207810 398792 214010 398848
rect 214066 398792 214071 398848
rect 207749 398790 214071 398792
rect 207749 398787 207815 398790
rect 214005 398787 214071 398790
rect 217182 398848 217291 398850
rect 217182 398792 217230 398848
rect 217286 398792 217291 398848
rect 217182 398787 217291 398792
rect 217501 398850 217567 398853
rect 217685 398850 217751 398853
rect 217501 398848 217751 398850
rect 217501 398792 217506 398848
rect 217562 398792 217690 398848
rect 217746 398792 217751 398848
rect 217501 398790 217751 398792
rect 217501 398787 217567 398790
rect 217685 398787 217751 398790
rect 216949 398714 217015 398717
rect 217182 398714 217242 398787
rect 216949 398712 217242 398714
rect 216949 398656 216954 398712
rect 217010 398656 217242 398712
rect 216949 398654 217242 398656
rect 219206 398714 219266 399062
rect 219341 399059 219407 399062
rect 229369 398986 229435 398989
rect 245377 398986 245443 398989
rect 229369 398984 229570 398986
rect 229369 398928 229374 398984
rect 229430 398928 229570 398984
rect 229369 398926 229570 398928
rect 229369 398923 229435 398926
rect 219341 398714 219407 398717
rect 219206 398712 219407 398714
rect 219206 398656 219346 398712
rect 219402 398656 219407 398712
rect 219206 398654 219407 398656
rect 216949 398651 217015 398654
rect 219341 398651 219407 398654
rect 211521 398578 211587 398581
rect 200070 398576 211587 398578
rect 200070 398520 211526 398576
rect 211582 398520 211587 398576
rect 200070 398518 211587 398520
rect 178677 398306 178743 398309
rect 200070 398306 200130 398518
rect 211521 398515 211587 398518
rect 202137 398442 202203 398445
rect 213361 398442 213427 398445
rect 202137 398440 213427 398442
rect 202137 398384 202142 398440
rect 202198 398384 213366 398440
rect 213422 398384 213427 398440
rect 202137 398382 213427 398384
rect 202137 398379 202203 398382
rect 213361 398379 213427 398382
rect 211153 398306 211219 398309
rect 178677 398304 200130 398306
rect 178677 398248 178682 398304
rect 178738 398248 200130 398304
rect 178677 398246 200130 398248
rect 209730 398304 211219 398306
rect 209730 398248 211158 398304
rect 211214 398248 211219 398304
rect 209730 398246 211219 398248
rect 178677 398243 178743 398246
rect 188337 398170 188403 398173
rect 209730 398170 209790 398246
rect 211153 398243 211219 398246
rect 212165 398306 212231 398309
rect 212441 398306 212507 398309
rect 212165 398304 212507 398306
rect 212165 398248 212170 398304
rect 212226 398248 212446 398304
rect 212502 398248 212507 398304
rect 212165 398246 212507 398248
rect 212165 398243 212231 398246
rect 212441 398243 212507 398246
rect 188337 398168 209790 398170
rect 188337 398112 188342 398168
rect 188398 398112 209790 398168
rect 188337 398110 209790 398112
rect 188337 398107 188403 398110
rect 228766 398108 228772 398172
rect 228836 398170 228842 398172
rect 229185 398170 229251 398173
rect 228836 398168 229251 398170
rect 228836 398112 229190 398168
rect 229246 398112 229251 398168
rect 228836 398110 229251 398112
rect 229510 398170 229570 398926
rect 245377 398984 253950 398986
rect 245377 398928 245382 398984
rect 245438 398928 253950 398984
rect 245377 398926 253950 398928
rect 245377 398923 245443 398926
rect 253890 398850 253950 398926
rect 302190 398926 314670 398986
rect 254526 398850 254532 398852
rect 253890 398790 254532 398850
rect 254526 398788 254532 398790
rect 254596 398788 254602 398852
rect 264278 398788 264284 398852
rect 264348 398850 264354 398852
rect 302190 398850 302250 398926
rect 264348 398790 302250 398850
rect 314610 398850 314670 398926
rect 337377 398850 337443 398853
rect 314610 398848 337443 398850
rect 314610 398792 337382 398848
rect 337438 398792 337443 398848
rect 314610 398790 337443 398792
rect 264348 398788 264354 398790
rect 337377 398787 337443 398790
rect 246481 398714 246547 398717
rect 246438 398712 246547 398714
rect 246438 398656 246486 398712
rect 246542 398656 246547 398712
rect 246438 398651 246547 398656
rect 248505 398714 248571 398717
rect 255957 398714 256023 398717
rect 248505 398712 256023 398714
rect 248505 398656 248510 398712
rect 248566 398656 255962 398712
rect 256018 398656 256023 398712
rect 248505 398654 256023 398656
rect 248505 398651 248571 398654
rect 255957 398651 256023 398654
rect 262806 398652 262812 398716
rect 262876 398714 262882 398716
rect 354121 398714 354187 398717
rect 262876 398712 354187 398714
rect 262876 398656 354126 398712
rect 354182 398656 354187 398712
rect 262876 398654 354187 398656
rect 262876 398652 262882 398654
rect 354121 398651 354187 398654
rect 246205 398306 246271 398309
rect 246438 398306 246498 398651
rect 247309 398578 247375 398581
rect 271137 398578 271203 398581
rect 247309 398576 271203 398578
rect 247309 398520 247314 398576
rect 247370 398520 271142 398576
rect 271198 398520 271203 398576
rect 247309 398518 271203 398520
rect 247309 398515 247375 398518
rect 271137 398515 271203 398518
rect 248505 398442 248571 398445
rect 249057 398442 249123 398445
rect 248505 398440 249123 398442
rect 248505 398384 248510 398440
rect 248566 398384 249062 398440
rect 249118 398384 249123 398440
rect 248505 398382 249123 398384
rect 248505 398379 248571 398382
rect 249057 398379 249123 398382
rect 255405 398442 255471 398445
rect 418797 398442 418863 398445
rect 255405 398440 418863 398442
rect 255405 398384 255410 398440
rect 255466 398384 418802 398440
rect 418858 398384 418863 398440
rect 255405 398382 418863 398384
rect 255405 398379 255471 398382
rect 418797 398379 418863 398382
rect 246205 398304 246498 398306
rect 246205 398248 246210 398304
rect 246266 398248 246498 398304
rect 246205 398246 246498 398248
rect 247309 398306 247375 398309
rect 247953 398306 248019 398309
rect 247309 398304 248019 398306
rect 247309 398248 247314 398304
rect 247370 398248 247958 398304
rect 248014 398248 248019 398304
rect 247309 398246 248019 398248
rect 246205 398243 246271 398246
rect 247309 398243 247375 398246
rect 247953 398243 248019 398246
rect 248781 398306 248847 398309
rect 494053 398306 494119 398309
rect 248781 398304 494119 398306
rect 248781 398248 248786 398304
rect 248842 398248 494058 398304
rect 494114 398248 494119 398304
rect 248781 398246 494119 398248
rect 248781 398243 248847 398246
rect 494053 398243 494119 398246
rect 229737 398170 229803 398173
rect 229510 398168 229803 398170
rect 229510 398112 229742 398168
rect 229798 398112 229803 398168
rect 229510 398110 229803 398112
rect 228836 398108 228842 398110
rect 229185 398107 229251 398110
rect 229737 398107 229803 398110
rect 242617 398170 242683 398173
rect 248781 398170 248847 398173
rect 242617 398168 248847 398170
rect 242617 398112 242622 398168
rect 242678 398112 248786 398168
rect 248842 398112 248847 398168
rect 242617 398110 248847 398112
rect 242617 398107 242683 398110
rect 248781 398107 248847 398110
rect 249885 398170 249951 398173
rect 507853 398170 507919 398173
rect 249885 398168 507919 398170
rect 249885 398112 249890 398168
rect 249946 398112 507858 398168
rect 507914 398112 507919 398168
rect 249885 398110 507919 398112
rect 249885 398107 249951 398110
rect 507853 398107 507919 398110
rect 25497 398034 25563 398037
rect 210693 398034 210759 398037
rect 212809 398034 212875 398037
rect 25497 398032 200130 398034
rect 25497 397976 25502 398032
rect 25558 397976 200130 398032
rect 25497 397974 200130 397976
rect 25497 397971 25563 397974
rect 200070 397898 200130 397974
rect 210693 398032 212875 398034
rect 210693 397976 210698 398032
rect 210754 397976 212814 398032
rect 212870 397976 212875 398032
rect 210693 397974 212875 397976
rect 210693 397971 210759 397974
rect 212809 397971 212875 397974
rect 251265 398034 251331 398037
rect 525793 398034 525859 398037
rect 251265 398032 525859 398034
rect 251265 397976 251270 398032
rect 251326 397976 525798 398032
rect 525854 397976 525859 398032
rect 251265 397974 525859 397976
rect 251265 397971 251331 397974
rect 525793 397971 525859 397974
rect 211889 397898 211955 397901
rect 200070 397896 211955 397898
rect 200070 397840 211894 397896
rect 211950 397840 211955 397896
rect 200070 397838 211955 397840
rect 211889 397835 211955 397838
rect 212257 397898 212323 397901
rect 215845 397898 215911 397901
rect 212257 397896 215911 397898
rect 212257 397840 212262 397896
rect 212318 397840 215850 397896
rect 215906 397840 215911 397896
rect 212257 397838 215911 397840
rect 212257 397835 212323 397838
rect 215845 397835 215911 397838
rect 216622 397836 216628 397900
rect 216692 397898 216698 397900
rect 217041 397898 217107 397901
rect 216692 397896 217107 397898
rect 216692 397840 217046 397896
rect 217102 397840 217107 397896
rect 216692 397838 217107 397840
rect 216692 397836 216698 397838
rect 217041 397835 217107 397838
rect 224953 397898 225019 397901
rect 225454 397898 225460 397900
rect 224953 397896 225460 397898
rect 224953 397840 224958 397896
rect 225014 397840 225460 397896
rect 224953 397838 225460 397840
rect 224953 397835 225019 397838
rect 225454 397836 225460 397838
rect 225524 397836 225530 397900
rect 230197 397898 230263 397901
rect 230422 397898 230428 397900
rect 230197 397896 230428 397898
rect 230197 397840 230202 397896
rect 230258 397840 230428 397896
rect 230197 397838 230428 397840
rect 230197 397835 230263 397838
rect 230422 397836 230428 397838
rect 230492 397836 230498 397900
rect 232957 397898 233023 397901
rect 233182 397898 233188 397900
rect 232957 397896 233188 397898
rect 232957 397840 232962 397896
rect 233018 397840 233188 397896
rect 232957 397838 233188 397840
rect 232957 397835 233023 397838
rect 233182 397836 233188 397838
rect 233252 397836 233258 397900
rect 242382 397836 242388 397900
rect 242452 397898 242458 397900
rect 242801 397898 242867 397901
rect 242452 397896 242867 397898
rect 242452 397840 242806 397896
rect 242862 397840 242867 397896
rect 242452 397838 242867 397840
rect 242452 397836 242458 397838
rect 242801 397835 242867 397838
rect 246757 397898 246823 397901
rect 246982 397898 246988 397900
rect 246757 397896 246988 397898
rect 246757 397840 246762 397896
rect 246818 397840 246988 397896
rect 246757 397838 246988 397840
rect 246757 397835 246823 397838
rect 246982 397836 246988 397838
rect 247052 397836 247058 397900
rect 247718 397836 247724 397900
rect 247788 397898 247794 397900
rect 248137 397898 248203 397901
rect 247788 397896 248203 397898
rect 247788 397840 248142 397896
rect 248198 397840 248203 397896
rect 247788 397838 248203 397840
rect 247788 397836 247794 397838
rect 248137 397835 248203 397838
rect 251950 397836 251956 397900
rect 252020 397898 252026 397900
rect 252461 397898 252527 397901
rect 252020 397896 252527 397898
rect 252020 397840 252466 397896
rect 252522 397840 252527 397896
rect 252020 397838 252527 397840
rect 252020 397836 252026 397838
rect 252461 397835 252527 397838
rect 254526 397836 254532 397900
rect 254596 397898 254602 397900
rect 260097 397898 260163 397901
rect 254596 397896 260163 397898
rect 254596 397840 260102 397896
rect 260158 397840 260163 397896
rect 254596 397838 260163 397840
rect 254596 397836 254602 397838
rect 260097 397835 260163 397838
rect 203609 397762 203675 397765
rect 210693 397762 210759 397765
rect 203609 397760 210759 397762
rect 203609 397704 203614 397760
rect 203670 397704 210698 397760
rect 210754 397704 210759 397760
rect 203609 397702 210759 397704
rect 203609 397699 203675 397702
rect 210693 397699 210759 397702
rect 211102 397700 211108 397764
rect 211172 397762 211178 397764
rect 211613 397762 211679 397765
rect 211172 397760 211679 397762
rect 211172 397704 211618 397760
rect 211674 397704 211679 397760
rect 211172 397702 211679 397704
rect 211172 397700 211178 397702
rect 211613 397699 211679 397702
rect 212533 397762 212599 397765
rect 212758 397762 212764 397764
rect 212533 397760 212764 397762
rect 212533 397704 212538 397760
rect 212594 397704 212764 397760
rect 212533 397702 212764 397704
rect 212533 397699 212599 397702
rect 212758 397700 212764 397702
rect 212828 397700 212834 397764
rect 214189 397762 214255 397765
rect 214414 397762 214420 397764
rect 214189 397760 214420 397762
rect 214189 397704 214194 397760
rect 214250 397704 214420 397760
rect 214189 397702 214420 397704
rect 214189 397699 214255 397702
rect 214414 397700 214420 397702
rect 214484 397700 214490 397764
rect 215334 397700 215340 397764
rect 215404 397762 215410 397764
rect 215569 397762 215635 397765
rect 215404 397760 215635 397762
rect 215404 397704 215574 397760
rect 215630 397704 215635 397760
rect 215404 397702 215635 397704
rect 215404 397700 215410 397702
rect 215569 397699 215635 397702
rect 216857 397762 216923 397765
rect 217174 397762 217180 397764
rect 216857 397760 217180 397762
rect 216857 397704 216862 397760
rect 216918 397704 217180 397760
rect 216857 397702 217180 397704
rect 216857 397699 216923 397702
rect 217174 397700 217180 397702
rect 217244 397700 217250 397764
rect 218237 397762 218303 397765
rect 219014 397762 219020 397764
rect 218237 397760 219020 397762
rect 218237 397704 218242 397760
rect 218298 397704 219020 397760
rect 218237 397702 219020 397704
rect 218237 397699 218303 397702
rect 219014 397700 219020 397702
rect 219084 397700 219090 397764
rect 220905 397762 220971 397765
rect 222193 397764 222259 397765
rect 221222 397762 221228 397764
rect 220905 397760 221228 397762
rect 220905 397704 220910 397760
rect 220966 397704 221228 397760
rect 220905 397702 221228 397704
rect 220905 397699 220971 397702
rect 221222 397700 221228 397702
rect 221292 397700 221298 397764
rect 222142 397762 222148 397764
rect 222102 397702 222148 397762
rect 222212 397760 222259 397764
rect 222254 397704 222259 397760
rect 222142 397700 222148 397702
rect 222212 397700 222259 397704
rect 222193 397699 222259 397700
rect 223573 397762 223639 397765
rect 223798 397762 223804 397764
rect 223573 397760 223804 397762
rect 223573 397704 223578 397760
rect 223634 397704 223804 397760
rect 223573 397702 223804 397704
rect 223573 397699 223639 397702
rect 223798 397700 223804 397702
rect 223868 397700 223874 397764
rect 224902 397700 224908 397764
rect 224972 397762 224978 397764
rect 225413 397762 225479 397765
rect 224972 397760 225479 397762
rect 224972 397704 225418 397760
rect 225474 397704 225479 397760
rect 224972 397702 225479 397704
rect 224972 397700 224978 397702
rect 225413 397699 225479 397702
rect 229870 397700 229876 397764
rect 229940 397762 229946 397764
rect 230381 397762 230447 397765
rect 229940 397760 230447 397762
rect 229940 397704 230386 397760
rect 230442 397704 230447 397760
rect 229940 397702 230447 397704
rect 229940 397700 229946 397702
rect 230381 397699 230447 397702
rect 230606 397700 230612 397764
rect 230676 397762 230682 397764
rect 231577 397762 231643 397765
rect 230676 397760 231643 397762
rect 230676 397704 231582 397760
rect 231638 397704 231643 397760
rect 230676 397702 231643 397704
rect 230676 397700 230682 397702
rect 231577 397699 231643 397702
rect 232630 397700 232636 397764
rect 232700 397762 232706 397764
rect 233141 397762 233207 397765
rect 232700 397760 233207 397762
rect 232700 397704 233146 397760
rect 233202 397704 233207 397760
rect 232700 397702 233207 397704
rect 232700 397700 232706 397702
rect 233141 397699 233207 397702
rect 233918 397700 233924 397764
rect 233988 397762 233994 397764
rect 234429 397762 234495 397765
rect 233988 397760 234495 397762
rect 233988 397704 234434 397760
rect 234490 397704 234495 397760
rect 233988 397702 234495 397704
rect 233988 397700 233994 397702
rect 234429 397699 234495 397702
rect 235206 397700 235212 397764
rect 235276 397762 235282 397764
rect 235901 397762 235967 397765
rect 235276 397760 235967 397762
rect 235276 397704 235906 397760
rect 235962 397704 235967 397760
rect 235276 397702 235967 397704
rect 235276 397700 235282 397702
rect 235901 397699 235967 397702
rect 236862 397700 236868 397764
rect 236932 397762 236938 397764
rect 237097 397762 237163 397765
rect 236932 397760 237163 397762
rect 236932 397704 237102 397760
rect 237158 397704 237163 397760
rect 236932 397702 237163 397704
rect 236932 397700 236938 397702
rect 237097 397699 237163 397702
rect 237966 397700 237972 397764
rect 238036 397762 238042 397764
rect 238569 397762 238635 397765
rect 238036 397760 238635 397762
rect 238036 397704 238574 397760
rect 238630 397704 238635 397760
rect 238036 397702 238635 397704
rect 238036 397700 238042 397702
rect 238569 397699 238635 397702
rect 239438 397700 239444 397764
rect 239508 397762 239514 397764
rect 240041 397762 240107 397765
rect 239508 397760 240107 397762
rect 239508 397704 240046 397760
rect 240102 397704 240107 397760
rect 239508 397702 240107 397704
rect 239508 397700 239514 397702
rect 240041 397699 240107 397702
rect 242198 397700 242204 397764
rect 242268 397762 242274 397764
rect 242525 397762 242591 397765
rect 242268 397760 242591 397762
rect 242268 397704 242530 397760
rect 242586 397704 242591 397760
rect 242268 397702 242591 397704
rect 242268 397700 242274 397702
rect 242525 397699 242591 397702
rect 243670 397700 243676 397764
rect 243740 397762 243746 397764
rect 244181 397762 244247 397765
rect 243740 397760 244247 397762
rect 243740 397704 244186 397760
rect 244242 397704 244247 397760
rect 243740 397702 244247 397704
rect 243740 397700 243746 397702
rect 244181 397699 244247 397702
rect 246614 397700 246620 397764
rect 246684 397762 246690 397764
rect 246941 397762 247007 397765
rect 246684 397760 247007 397762
rect 246684 397704 246946 397760
rect 247002 397704 247007 397760
rect 246684 397702 247007 397704
rect 246684 397700 246690 397702
rect 246941 397699 247007 397702
rect 247902 397700 247908 397764
rect 247972 397762 247978 397764
rect 248229 397762 248295 397765
rect 247972 397760 248295 397762
rect 247972 397704 248234 397760
rect 248290 397704 248295 397760
rect 247972 397702 248295 397704
rect 247972 397700 247978 397702
rect 248229 397699 248295 397702
rect 248638 397700 248644 397764
rect 248708 397762 248714 397764
rect 249701 397762 249767 397765
rect 248708 397760 249767 397762
rect 248708 397704 249706 397760
rect 249762 397704 249767 397760
rect 248708 397702 249767 397704
rect 248708 397700 248714 397702
rect 249701 397699 249767 397702
rect 250662 397700 250668 397764
rect 250732 397762 250738 397764
rect 251081 397762 251147 397765
rect 250732 397760 251147 397762
rect 250732 397704 251086 397760
rect 251142 397704 251147 397760
rect 250732 397702 251147 397704
rect 250732 397700 250738 397702
rect 251081 397699 251147 397702
rect 251766 397700 251772 397764
rect 251836 397762 251842 397764
rect 252185 397762 252251 397765
rect 251836 397760 252251 397762
rect 251836 397704 252190 397760
rect 252246 397704 252251 397760
rect 251836 397702 252251 397704
rect 251836 397700 251842 397702
rect 252185 397699 252251 397702
rect 253422 397700 253428 397764
rect 253492 397762 253498 397764
rect 253841 397762 253907 397765
rect 253492 397760 253907 397762
rect 253492 397704 253846 397760
rect 253902 397704 253907 397760
rect 253492 397702 253907 397704
rect 253492 397700 253498 397702
rect 253841 397699 253907 397702
rect 254710 397700 254716 397764
rect 254780 397762 254786 397764
rect 255221 397762 255287 397765
rect 254780 397760 255287 397762
rect 254780 397704 255226 397760
rect 255282 397704 255287 397760
rect 254780 397702 255287 397704
rect 254780 397700 254786 397702
rect 255221 397699 255287 397702
rect 211429 397628 211495 397629
rect 211429 397624 211476 397628
rect 211540 397626 211546 397628
rect 211797 397626 211863 397629
rect 212993 397626 213059 397629
rect -960 397490 480 397580
rect 211429 397568 211434 397624
rect 211429 397564 211476 397568
rect 211540 397566 211586 397626
rect 211797 397624 213059 397626
rect 211797 397568 211802 397624
rect 211858 397568 212998 397624
rect 213054 397568 213059 397624
rect 211797 397566 213059 397568
rect 211540 397564 211546 397566
rect 211429 397563 211495 397564
rect 211797 397563 211863 397566
rect 212993 397563 213059 397566
rect 214046 397564 214052 397628
rect 214116 397626 214122 397628
rect 214281 397626 214347 397629
rect 214116 397624 214347 397626
rect 214116 397568 214286 397624
rect 214342 397568 214347 397624
rect 214116 397566 214347 397568
rect 214116 397564 214122 397566
rect 214281 397563 214347 397566
rect 215477 397626 215543 397629
rect 215702 397626 215708 397628
rect 215477 397624 215708 397626
rect 215477 397568 215482 397624
rect 215538 397568 215708 397624
rect 215477 397566 215708 397568
rect 215477 397563 215543 397566
rect 215702 397564 215708 397566
rect 215772 397564 215778 397628
rect 216673 397626 216739 397629
rect 216990 397626 216996 397628
rect 216673 397624 216996 397626
rect 216673 397568 216678 397624
rect 216734 397568 216996 397624
rect 216673 397566 216996 397568
rect 216673 397563 216739 397566
rect 216990 397564 216996 397566
rect 217060 397564 217066 397628
rect 218053 397626 218119 397629
rect 218830 397626 218836 397628
rect 218053 397624 218836 397626
rect 218053 397568 218058 397624
rect 218114 397568 218836 397624
rect 218053 397566 218836 397568
rect 218053 397563 218119 397566
rect 218830 397564 218836 397566
rect 218900 397564 218906 397628
rect 219566 397564 219572 397628
rect 219636 397626 219642 397628
rect 219801 397626 219867 397629
rect 219636 397624 219867 397626
rect 219636 397568 219806 397624
rect 219862 397568 219867 397624
rect 219636 397566 219867 397568
rect 219636 397564 219642 397566
rect 219801 397563 219867 397566
rect 220854 397564 220860 397628
rect 220924 397626 220930 397628
rect 220997 397626 221063 397629
rect 220924 397624 221063 397626
rect 220924 397568 221002 397624
rect 221058 397568 221063 397624
rect 220924 397566 221063 397568
rect 220924 397564 220930 397566
rect 220997 397563 221063 397566
rect 221181 397626 221247 397629
rect 221406 397626 221412 397628
rect 221181 397624 221412 397626
rect 221181 397568 221186 397624
rect 221242 397568 221412 397624
rect 221181 397566 221412 397568
rect 221181 397563 221247 397566
rect 221406 397564 221412 397566
rect 221476 397564 221482 397628
rect 223849 397626 223915 397629
rect 225137 397628 225203 397629
rect 223982 397626 223988 397628
rect 223849 397624 223988 397626
rect 223849 397568 223854 397624
rect 223910 397568 223988 397624
rect 223849 397566 223988 397568
rect 223849 397563 223915 397566
rect 223982 397564 223988 397566
rect 224052 397564 224058 397628
rect 225086 397626 225092 397628
rect 225046 397566 225092 397626
rect 225156 397624 225203 397628
rect 225198 397568 225203 397624
rect 225086 397564 225092 397566
rect 225156 397564 225203 397568
rect 225137 397563 225203 397564
rect 226517 397628 226583 397629
rect 226517 397624 226564 397628
rect 226628 397626 226634 397628
rect 226517 397568 226522 397624
rect 226517 397564 226564 397568
rect 226628 397566 226674 397626
rect 226628 397564 226634 397566
rect 228582 397564 228588 397628
rect 228652 397626 228658 397628
rect 229001 397626 229067 397629
rect 230105 397628 230171 397629
rect 230054 397626 230060 397628
rect 228652 397624 229067 397626
rect 228652 397568 229006 397624
rect 229062 397568 229067 397624
rect 228652 397566 229067 397568
rect 230014 397566 230060 397626
rect 230124 397624 230171 397628
rect 230166 397568 230171 397624
rect 228652 397564 228658 397566
rect 226517 397563 226583 397564
rect 229001 397563 229067 397566
rect 230054 397564 230060 397566
rect 230124 397564 230171 397568
rect 230790 397564 230796 397628
rect 230860 397626 230866 397628
rect 231761 397626 231827 397629
rect 232865 397628 232931 397629
rect 232814 397626 232820 397628
rect 230860 397624 231827 397626
rect 230860 397568 231766 397624
rect 231822 397568 231827 397624
rect 230860 397566 231827 397568
rect 232774 397566 232820 397626
rect 232884 397624 232931 397628
rect 232926 397568 232931 397624
rect 230860 397564 230866 397566
rect 230105 397563 230171 397564
rect 231761 397563 231827 397566
rect 232814 397564 232820 397566
rect 232884 397564 232931 397568
rect 234102 397564 234108 397628
rect 234172 397626 234178 397628
rect 234337 397626 234403 397629
rect 234172 397624 234403 397626
rect 234172 397568 234342 397624
rect 234398 397568 234403 397624
rect 234172 397566 234403 397568
rect 234172 397564 234178 397566
rect 232865 397563 232931 397564
rect 234337 397563 234403 397566
rect 235390 397564 235396 397628
rect 235460 397626 235466 397628
rect 235717 397626 235783 397629
rect 235460 397624 235783 397626
rect 235460 397568 235722 397624
rect 235778 397568 235783 397624
rect 235460 397566 235783 397568
rect 235460 397564 235466 397566
rect 235717 397563 235783 397566
rect 237046 397564 237052 397628
rect 237116 397626 237122 397628
rect 237281 397626 237347 397629
rect 237116 397624 237347 397626
rect 237116 397568 237286 397624
rect 237342 397568 237347 397624
rect 237116 397566 237347 397568
rect 237116 397564 237122 397566
rect 237281 397563 237347 397566
rect 238150 397564 238156 397628
rect 238220 397626 238226 397628
rect 238477 397626 238543 397629
rect 238220 397624 238543 397626
rect 238220 397568 238482 397624
rect 238538 397568 238543 397624
rect 238220 397566 238543 397568
rect 238220 397564 238226 397566
rect 238477 397563 238543 397566
rect 239622 397564 239628 397628
rect 239692 397626 239698 397628
rect 239765 397626 239831 397629
rect 239692 397624 239831 397626
rect 239692 397568 239770 397624
rect 239826 397568 239831 397624
rect 239692 397566 239831 397568
rect 239692 397564 239698 397566
rect 239765 397563 239831 397566
rect 242433 397626 242499 397629
rect 242750 397626 242756 397628
rect 242433 397624 242756 397626
rect 242433 397568 242438 397624
rect 242494 397568 242756 397624
rect 242433 397566 242756 397568
rect 242433 397563 242499 397566
rect 242750 397564 242756 397566
rect 242820 397564 242826 397628
rect 243854 397564 243860 397628
rect 243924 397626 243930 397628
rect 243997 397626 244063 397629
rect 243924 397624 244063 397626
rect 243924 397568 244002 397624
rect 244058 397568 244063 397624
rect 243924 397566 244063 397568
rect 243924 397564 243930 397566
rect 243997 397563 244063 397566
rect 246430 397564 246436 397628
rect 246500 397626 246506 397628
rect 246665 397626 246731 397629
rect 246500 397624 246731 397626
rect 246500 397568 246670 397624
rect 246726 397568 246731 397624
rect 246500 397566 246731 397568
rect 246500 397564 246506 397566
rect 246665 397563 246731 397566
rect 248086 397564 248092 397628
rect 248156 397626 248162 397628
rect 248321 397626 248387 397629
rect 248156 397624 248387 397626
rect 248156 397568 248326 397624
rect 248382 397568 248387 397624
rect 248156 397566 248387 397568
rect 248156 397564 248162 397566
rect 248321 397563 248387 397566
rect 248822 397564 248828 397628
rect 248892 397626 248898 397628
rect 249517 397626 249583 397629
rect 250805 397628 250871 397629
rect 250805 397626 250852 397628
rect 248892 397624 249583 397626
rect 248892 397568 249522 397624
rect 249578 397568 249583 397624
rect 248892 397566 249583 397568
rect 250760 397624 250852 397626
rect 250760 397568 250810 397624
rect 250760 397566 250852 397568
rect 248892 397564 248898 397566
rect 249517 397563 249583 397566
rect 250805 397564 250852 397566
rect 250916 397564 250922 397628
rect 252134 397564 252140 397628
rect 252204 397626 252210 397628
rect 252277 397626 252343 397629
rect 252204 397624 252343 397626
rect 252204 397568 252282 397624
rect 252338 397568 252343 397624
rect 252204 397566 252343 397568
rect 252204 397564 252210 397566
rect 250805 397563 250871 397564
rect 252277 397563 252343 397566
rect 253238 397564 253244 397628
rect 253308 397626 253314 397628
rect 253565 397626 253631 397629
rect 253308 397624 253631 397626
rect 253308 397568 253570 397624
rect 253626 397568 253631 397624
rect 253308 397566 253631 397568
rect 253308 397564 253314 397566
rect 253565 397563 253631 397566
rect 254894 397564 254900 397628
rect 254964 397626 254970 397628
rect 255037 397626 255103 397629
rect 254964 397624 255103 397626
rect 254964 397568 255042 397624
rect 255098 397568 255103 397624
rect 254964 397566 255103 397568
rect 254964 397564 254970 397566
rect 255037 397563 255103 397566
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 209814 397428 209820 397492
rect 209884 397490 209890 397492
rect 210325 397490 210391 397493
rect 211337 397492 211403 397493
rect 212625 397492 212691 397493
rect 211286 397490 211292 397492
rect 209884 397488 210391 397490
rect 209884 397432 210330 397488
rect 210386 397432 210391 397488
rect 209884 397430 210391 397432
rect 211246 397430 211292 397490
rect 211356 397488 211403 397492
rect 212574 397490 212580 397492
rect 211398 397432 211403 397488
rect 209884 397428 209890 397430
rect 210325 397427 210391 397430
rect 211286 397428 211292 397430
rect 211356 397428 211403 397432
rect 212534 397430 212580 397490
rect 212644 397488 212691 397492
rect 212686 397432 212691 397488
rect 212574 397428 212580 397430
rect 212644 397428 212691 397432
rect 211337 397427 211403 397428
rect 212625 397427 212691 397428
rect 214097 397490 214163 397493
rect 214230 397490 214236 397492
rect 214097 397488 214236 397490
rect 214097 397432 214102 397488
rect 214158 397432 214236 397488
rect 214097 397430 214236 397432
rect 214097 397427 214163 397430
rect 214230 397428 214236 397430
rect 214300 397428 214306 397492
rect 215293 397490 215359 397493
rect 216765 397492 216831 397493
rect 215518 397490 215524 397492
rect 215293 397488 215524 397490
rect 215293 397432 215298 397488
rect 215354 397432 215524 397488
rect 215293 397430 215524 397432
rect 215293 397427 215359 397430
rect 215518 397428 215524 397430
rect 215588 397428 215594 397492
rect 216765 397490 216812 397492
rect 216720 397488 216812 397490
rect 216720 397432 216770 397488
rect 216720 397430 216812 397432
rect 216765 397428 216812 397430
rect 216876 397428 216882 397492
rect 218145 397490 218211 397493
rect 218646 397490 218652 397492
rect 218145 397488 218652 397490
rect 218145 397432 218150 397488
rect 218206 397432 218652 397488
rect 218145 397430 218652 397432
rect 216765 397427 216831 397428
rect 218145 397427 218211 397430
rect 218646 397428 218652 397430
rect 218716 397428 218722 397492
rect 219382 397428 219388 397492
rect 219452 397490 219458 397492
rect 219525 397490 219591 397493
rect 219709 397492 219775 397493
rect 221089 397492 221155 397493
rect 219709 397490 219756 397492
rect 219452 397488 219591 397490
rect 219452 397432 219530 397488
rect 219586 397432 219591 397488
rect 219452 397430 219591 397432
rect 219664 397488 219756 397490
rect 219664 397432 219714 397488
rect 219664 397430 219756 397432
rect 219452 397428 219458 397430
rect 219525 397427 219591 397430
rect 219709 397428 219756 397430
rect 219820 397428 219826 397492
rect 221038 397490 221044 397492
rect 220998 397430 221044 397490
rect 221108 397488 221155 397492
rect 221150 397432 221155 397488
rect 221038 397428 221044 397430
rect 221108 397428 221155 397432
rect 219709 397427 219775 397428
rect 221089 397427 221155 397428
rect 222285 397490 222351 397493
rect 223062 397490 223068 397492
rect 222285 397488 223068 397490
rect 222285 397432 222290 397488
rect 222346 397432 223068 397488
rect 222285 397430 223068 397432
rect 222285 397427 222351 397430
rect 223062 397428 223068 397430
rect 223132 397428 223138 397492
rect 223614 397428 223620 397492
rect 223684 397490 223690 397492
rect 223757 397490 223823 397493
rect 223684 397488 223823 397490
rect 223684 397432 223762 397488
rect 223818 397432 223823 397488
rect 223684 397430 223823 397432
rect 223684 397428 223690 397430
rect 223757 397427 223823 397430
rect 223941 397490 224007 397493
rect 225229 397492 225295 397493
rect 226333 397492 226399 397493
rect 228909 397492 228975 397493
rect 230289 397492 230355 397493
rect 224166 397490 224172 397492
rect 223941 397488 224172 397490
rect 223941 397432 223946 397488
rect 224002 397432 224172 397488
rect 223941 397430 224172 397432
rect 223941 397427 224007 397430
rect 224166 397428 224172 397430
rect 224236 397428 224242 397492
rect 225229 397488 225276 397492
rect 225340 397490 225346 397492
rect 225229 397432 225234 397488
rect 225229 397428 225276 397432
rect 225340 397430 225386 397490
rect 226333 397488 226380 397492
rect 226444 397490 226450 397492
rect 226333 397432 226338 397488
rect 225340 397428 225346 397430
rect 226333 397428 226380 397432
rect 226444 397430 226490 397490
rect 228909 397488 228956 397492
rect 229020 397490 229026 397492
rect 230238 397490 230244 397492
rect 228909 397432 228914 397488
rect 226444 397428 226450 397430
rect 228909 397428 228956 397432
rect 229020 397430 229066 397490
rect 230198 397430 230244 397490
rect 230308 397488 230355 397492
rect 230350 397432 230355 397488
rect 229020 397428 229026 397430
rect 230238 397428 230244 397430
rect 230308 397428 230355 397432
rect 230974 397428 230980 397492
rect 231044 397490 231050 397492
rect 231669 397490 231735 397493
rect 233049 397492 233115 397493
rect 232998 397490 233004 397492
rect 231044 397488 231735 397490
rect 231044 397432 231674 397488
rect 231730 397432 231735 397488
rect 231044 397430 231735 397432
rect 232958 397430 233004 397490
rect 233068 397488 233115 397492
rect 233110 397432 233115 397488
rect 231044 397428 231050 397430
rect 225229 397427 225295 397428
rect 226333 397427 226399 397428
rect 228909 397427 228975 397428
rect 230289 397427 230355 397428
rect 231669 397427 231735 397430
rect 232998 397428 233004 397430
rect 233068 397428 233115 397432
rect 233049 397427 233115 397428
rect 234245 397492 234311 397493
rect 234245 397488 234292 397492
rect 234356 397490 234362 397492
rect 234245 397432 234250 397488
rect 234245 397428 234292 397432
rect 234356 397430 234402 397490
rect 234356 397428 234362 397430
rect 235574 397428 235580 397492
rect 235644 397490 235650 397492
rect 235809 397490 235875 397493
rect 235644 397488 235875 397490
rect 235644 397432 235814 397488
rect 235870 397432 235875 397488
rect 235644 397430 235875 397432
rect 235644 397428 235650 397430
rect 234245 397427 234311 397428
rect 235809 397427 235875 397430
rect 237189 397492 237255 397493
rect 238385 397492 238451 397493
rect 237189 397488 237236 397492
rect 237300 397490 237306 397492
rect 238334 397490 238340 397492
rect 237189 397432 237194 397488
rect 237189 397428 237236 397432
rect 237300 397430 237346 397490
rect 238294 397430 238340 397490
rect 238404 397488 238451 397492
rect 238446 397432 238451 397488
rect 237300 397428 237306 397430
rect 238334 397428 238340 397430
rect 238404 397428 238451 397432
rect 237189 397427 237255 397428
rect 238385 397427 238451 397428
rect 239673 397490 239739 397493
rect 239949 397492 240015 397493
rect 239806 397490 239812 397492
rect 239673 397488 239812 397490
rect 239673 397432 239678 397488
rect 239734 397432 239812 397488
rect 239673 397430 239812 397432
rect 239673 397427 239739 397430
rect 239806 397428 239812 397430
rect 239876 397428 239882 397492
rect 239949 397488 239996 397492
rect 240060 397490 240066 397492
rect 239949 397432 239954 397488
rect 239949 397428 239996 397432
rect 240060 397430 240106 397490
rect 240060 397428 240066 397430
rect 241094 397428 241100 397492
rect 241164 397490 241170 397492
rect 241329 397490 241395 397493
rect 241164 397488 241395 397490
rect 241164 397432 241334 397488
rect 241390 397432 241395 397488
rect 241164 397430 241395 397432
rect 241164 397428 241170 397430
rect 239949 397427 240015 397428
rect 241329 397427 241395 397430
rect 242566 397428 242572 397492
rect 242636 397490 242642 397492
rect 242709 397490 242775 397493
rect 244089 397492 244155 397493
rect 244038 397490 244044 397492
rect 242636 397488 242775 397490
rect 242636 397432 242714 397488
rect 242770 397432 242775 397488
rect 242636 397430 242775 397432
rect 243998 397430 244044 397490
rect 244108 397488 244155 397492
rect 245469 397492 245535 397493
rect 246849 397492 246915 397493
rect 245469 397490 245516 397492
rect 244150 397432 244155 397488
rect 242636 397428 242642 397430
rect 242709 397427 242775 397430
rect 244038 397428 244044 397430
rect 244108 397428 244155 397432
rect 245424 397488 245516 397490
rect 245424 397432 245474 397488
rect 245424 397430 245516 397432
rect 244089 397427 244155 397428
rect 245469 397428 245516 397430
rect 245580 397428 245586 397492
rect 246798 397490 246804 397492
rect 246758 397430 246804 397490
rect 246868 397488 246915 397492
rect 246910 397432 246915 397488
rect 246798 397428 246804 397430
rect 246868 397428 246915 397432
rect 245469 397427 245535 397428
rect 246849 397427 246915 397428
rect 248045 397490 248111 397493
rect 248270 397490 248276 397492
rect 248045 397488 248276 397490
rect 248045 397432 248050 397488
rect 248106 397432 248276 397488
rect 248045 397430 248276 397432
rect 248045 397427 248111 397430
rect 248270 397428 248276 397430
rect 248340 397428 248346 397492
rect 249006 397428 249012 397492
rect 249076 397490 249082 397492
rect 249609 397490 249675 397493
rect 250989 397492 251055 397493
rect 252369 397492 252435 397493
rect 250989 397490 251036 397492
rect 249076 397488 249675 397490
rect 249076 397432 249614 397488
rect 249670 397432 249675 397488
rect 249076 397430 249675 397432
rect 250944 397488 251036 397490
rect 250944 397432 250994 397488
rect 250944 397430 251036 397432
rect 249076 397428 249082 397430
rect 249609 397427 249675 397430
rect 250989 397428 251036 397430
rect 251100 397428 251106 397492
rect 252318 397490 252324 397492
rect 252278 397430 252324 397490
rect 252388 397488 252435 397492
rect 252430 397432 252435 397488
rect 252318 397428 252324 397430
rect 252388 397428 252435 397432
rect 253606 397428 253612 397492
rect 253676 397490 253682 397492
rect 253749 397490 253815 397493
rect 255129 397492 255195 397493
rect 255078 397490 255084 397492
rect 253676 397488 253815 397490
rect 253676 397432 253754 397488
rect 253810 397432 253815 397488
rect 253676 397430 253815 397432
rect 255038 397430 255084 397490
rect 255148 397488 255195 397492
rect 255190 397432 255195 397488
rect 253676 397428 253682 397430
rect 250989 397427 251055 397428
rect 252369 397427 252435 397428
rect 253749 397427 253815 397430
rect 255078 397428 255084 397430
rect 255148 397428 255195 397432
rect 255129 397427 255195 397428
rect 235625 397354 235691 397357
rect 324313 397354 324379 397357
rect 235625 397352 324379 397354
rect 235625 397296 235630 397352
rect 235686 397296 324318 397352
rect 324374 397296 324379 397352
rect 235625 397294 324379 397296
rect 235625 397291 235691 397294
rect 324313 397291 324379 397294
rect 238661 397218 238727 397221
rect 364333 397218 364399 397221
rect 238661 397216 364399 397218
rect 238661 397160 238666 397216
rect 238722 397160 364338 397216
rect 364394 397160 364399 397216
rect 238661 397158 364399 397160
rect 238661 397155 238727 397158
rect 364333 397155 364399 397158
rect 210325 397082 210391 397085
rect 215385 397082 215451 397085
rect 210325 397080 215451 397082
rect 210325 397024 210330 397080
rect 210386 397024 215390 397080
rect 215446 397024 215451 397080
rect 210325 397022 215451 397024
rect 210325 397019 210391 397022
rect 215385 397019 215451 397022
rect 241421 397082 241487 397085
rect 247033 397082 247099 397085
rect 398833 397082 398899 397085
rect 241421 397080 243738 397082
rect 241421 397024 241426 397080
rect 241482 397024 243738 397080
rect 241421 397022 243738 397024
rect 241421 397019 241487 397022
rect 151813 396946 151879 396949
rect 222142 396946 222148 396948
rect 151813 396944 222148 396946
rect 151813 396888 151818 396944
rect 151874 396888 222148 396944
rect 151813 396886 222148 396888
rect 151813 396883 151879 396886
rect 222142 396884 222148 396886
rect 222212 396884 222218 396948
rect 64873 396810 64939 396813
rect 210325 396810 210391 396813
rect 211245 396810 211311 396813
rect 232589 396810 232655 396813
rect 64873 396808 210391 396810
rect 64873 396752 64878 396808
rect 64934 396752 210330 396808
rect 210386 396752 210391 396808
rect 64873 396750 210391 396752
rect 64873 396747 64939 396750
rect 210325 396747 210391 396750
rect 210558 396808 211311 396810
rect 210558 396752 211250 396808
rect 211306 396752 211311 396808
rect 210558 396750 211311 396752
rect 11053 396674 11119 396677
rect 210558 396674 210618 396750
rect 211245 396747 211311 396750
rect 232454 396808 232655 396810
rect 232454 396752 232594 396808
rect 232650 396752 232655 396808
rect 232454 396750 232655 396752
rect 11053 396672 210618 396674
rect 11053 396616 11058 396672
rect 11114 396616 210618 396672
rect 11053 396614 210618 396616
rect 11053 396611 11119 396614
rect 232129 396538 232195 396541
rect 232454 396538 232514 396750
rect 232589 396747 232655 396750
rect 238845 396810 238911 396813
rect 239121 396810 239187 396813
rect 238845 396808 239187 396810
rect 238845 396752 238850 396808
rect 238906 396752 239126 396808
rect 239182 396752 239187 396808
rect 238845 396750 239187 396752
rect 238845 396747 238911 396750
rect 239121 396747 239187 396750
rect 243678 396674 243738 397022
rect 247033 397080 398899 397082
rect 247033 397024 247038 397080
rect 247094 397024 398838 397080
rect 398894 397024 398899 397080
rect 247033 397022 398899 397024
rect 247033 397019 247099 397022
rect 398833 397019 398899 397022
rect 243905 396946 243971 396949
rect 431953 396946 432019 396949
rect 243905 396944 432019 396946
rect 243905 396888 243910 396944
rect 243966 396888 431958 396944
rect 432014 396888 432019 396944
rect 243905 396886 432019 396888
rect 243905 396883 243971 396886
rect 431953 396883 432019 396886
rect 245561 396810 245627 396813
rect 452653 396810 452719 396813
rect 245561 396808 452719 396810
rect 245561 396752 245566 396808
rect 245622 396752 452658 396808
rect 452714 396752 452719 396808
rect 245561 396750 452719 396752
rect 245561 396747 245627 396750
rect 452653 396747 452719 396750
rect 247033 396674 247099 396677
rect 243678 396672 247099 396674
rect 243678 396616 247038 396672
rect 247094 396616 247099 396672
rect 243678 396614 247099 396616
rect 247033 396611 247099 396614
rect 250897 396674 250963 396677
rect 521653 396674 521719 396677
rect 250897 396672 521719 396674
rect 250897 396616 250902 396672
rect 250958 396616 521658 396672
rect 521714 396616 521719 396672
rect 250897 396614 521719 396616
rect 250897 396611 250963 396614
rect 521653 396611 521719 396614
rect 232129 396536 232514 396538
rect 232129 396480 232134 396536
rect 232190 396480 232514 396536
rect 232129 396478 232514 396480
rect 234429 396538 234495 396541
rect 310513 396538 310579 396541
rect 234429 396536 310579 396538
rect 234429 396480 234434 396536
rect 234490 396480 310518 396536
rect 310574 396480 310579 396536
rect 234429 396478 310579 396480
rect 232129 396475 232195 396478
rect 234429 396475 234495 396478
rect 310513 396475 310579 396478
rect 118693 395722 118759 395725
rect 219617 395722 219683 395725
rect 118693 395720 219683 395722
rect 118693 395664 118698 395720
rect 118754 395664 219622 395720
rect 219678 395664 219683 395720
rect 118693 395662 219683 395664
rect 118693 395659 118759 395662
rect 219617 395659 219683 395662
rect 67633 395586 67699 395589
rect 215334 395586 215340 395588
rect 67633 395584 215340 395586
rect 67633 395528 67638 395584
rect 67694 395528 215340 395584
rect 67633 395526 215340 395528
rect 67633 395523 67699 395526
rect 215334 395524 215340 395526
rect 215404 395524 215410 395588
rect 246982 395524 246988 395588
rect 247052 395586 247058 395588
rect 257337 395586 257403 395589
rect 247052 395584 257403 395586
rect 247052 395528 257342 395584
rect 257398 395528 257403 395584
rect 247052 395526 257403 395528
rect 247052 395524 247058 395526
rect 257337 395523 257403 395526
rect 45553 395450 45619 395453
rect 213913 395450 213979 395453
rect 45553 395448 213979 395450
rect 45553 395392 45558 395448
rect 45614 395392 213918 395448
rect 213974 395392 213979 395448
rect 45553 395390 213979 395392
rect 45553 395387 45619 395390
rect 213913 395387 213979 395390
rect 230422 395388 230428 395452
rect 230492 395450 230498 395452
rect 255221 395450 255287 395453
rect 230492 395448 255287 395450
rect 230492 395392 255226 395448
rect 255282 395392 255287 395448
rect 230492 395390 255287 395392
rect 230492 395388 230498 395390
rect 255221 395387 255287 395390
rect 27705 395314 27771 395317
rect 212758 395314 212764 395316
rect 27705 395312 212764 395314
rect 27705 395256 27710 395312
rect 27766 395256 212764 395312
rect 27705 395254 212764 395256
rect 27705 395251 27771 395254
rect 212758 395252 212764 395254
rect 212828 395252 212834 395316
rect 253054 395252 253060 395316
rect 253124 395314 253130 395316
rect 556153 395314 556219 395317
rect 253124 395312 556219 395314
rect 253124 395256 556158 395312
rect 556214 395256 556219 395312
rect 253124 395254 556219 395256
rect 253124 395252 253130 395254
rect 556153 395251 556219 395254
rect 213269 394770 213335 394773
rect 221222 394770 221228 394772
rect 213269 394768 221228 394770
rect 213269 394712 213274 394768
rect 213330 394712 221228 394768
rect 213269 394710 221228 394712
rect 213269 394707 213335 394710
rect 221222 394708 221228 394710
rect 221292 394708 221298 394772
rect 139393 393954 139459 393957
rect 221406 393954 221412 393956
rect 139393 393952 221412 393954
rect 139393 393896 139398 393952
rect 139454 393896 221412 393952
rect 139393 393894 221412 393896
rect 139393 393891 139459 393894
rect 221406 393892 221412 393894
rect 221476 393892 221482 393956
rect 233182 393892 233188 393956
rect 233252 393954 233258 393956
rect 291193 393954 291259 393957
rect 233252 393952 291259 393954
rect 233252 393896 291198 393952
rect 291254 393896 291259 393952
rect 233252 393894 291259 393896
rect 233252 393892 233258 393894
rect 291193 393891 291259 393894
rect 215937 393818 216003 393821
rect 215894 393816 216003 393818
rect 215894 393760 215942 393816
rect 215998 393760 216003 393816
rect 215894 393755 216003 393760
rect 215753 393546 215819 393549
rect 215894 393546 215954 393755
rect 215753 393544 215954 393546
rect 215753 393488 215758 393544
rect 215814 393488 215954 393544
rect 215753 393486 215954 393488
rect 215753 393483 215819 393486
rect 208393 392866 208459 392869
rect 226558 392866 226564 392868
rect 208393 392864 226564 392866
rect 208393 392808 208398 392864
rect 208454 392808 226564 392864
rect 208393 392806 226564 392808
rect 208393 392803 208459 392806
rect 226558 392804 226564 392806
rect 226628 392804 226634 392868
rect 187693 392730 187759 392733
rect 225454 392730 225460 392732
rect 187693 392728 225460 392730
rect 187693 392672 187698 392728
rect 187754 392672 225460 392728
rect 187693 392670 225460 392672
rect 187693 392667 187759 392670
rect 225454 392668 225460 392670
rect 225524 392668 225530 392732
rect 28993 392594 29059 392597
rect 212574 392594 212580 392596
rect 28993 392592 212580 392594
rect 28993 392536 28998 392592
rect 29054 392536 212580 392592
rect 28993 392534 212580 392536
rect 28993 392531 29059 392534
rect 212574 392532 212580 392534
rect 212644 392532 212650 392596
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 102133 355330 102199 355333
rect 219014 355330 219020 355332
rect 102133 355328 219020 355330
rect 102133 355272 102138 355328
rect 102194 355272 219020 355328
rect 102133 355270 219020 355272
rect 102133 355267 102199 355270
rect 219014 355268 219020 355270
rect 219084 355268 219090 355332
rect 235206 355268 235212 355332
rect 235276 355330 235282 355332
rect 328453 355330 328519 355333
rect 235276 355328 328519 355330
rect 235276 355272 328458 355328
rect 328514 355272 328519 355328
rect 235276 355270 328519 355272
rect 235276 355268 235282 355270
rect 328453 355267 328519 355270
rect 238150 354044 238156 354108
rect 238220 354106 238226 354108
rect 361573 354106 361639 354109
rect 238220 354104 361639 354106
rect 238220 354048 361578 354104
rect 361634 354048 361639 354104
rect 238220 354046 361639 354048
rect 238220 354044 238226 354046
rect 361573 354043 361639 354046
rect 251766 353908 251772 353972
rect 251836 353970 251842 353972
rect 538213 353970 538279 353973
rect 251836 353968 538279 353970
rect 251836 353912 538218 353968
rect 538274 353912 538279 353968
rect 251836 353910 538279 353912
rect 251836 353908 251842 353910
rect 538213 353907 538279 353910
rect 243670 352820 243676 352884
rect 243740 352882 243746 352884
rect 434713 352882 434779 352885
rect 243740 352880 434779 352882
rect 243740 352824 434718 352880
rect 434774 352824 434779 352880
rect 243740 352822 434779 352824
rect 243740 352820 243746 352822
rect 434713 352819 434779 352822
rect 247718 352684 247724 352748
rect 247788 352746 247794 352748
rect 485773 352746 485839 352749
rect 247788 352744 485839 352746
rect 247788 352688 485778 352744
rect 485834 352688 485839 352744
rect 247788 352686 485839 352688
rect 247788 352684 247794 352686
rect 485773 352683 485839 352686
rect 153193 352610 153259 352613
rect 223062 352610 223068 352612
rect 153193 352608 223068 352610
rect 153193 352552 153198 352608
rect 153254 352552 223068 352608
rect 153193 352550 223068 352552
rect 153193 352547 153259 352550
rect 223062 352548 223068 352550
rect 223132 352548 223138 352612
rect 248638 352548 248644 352612
rect 248708 352610 248714 352612
rect 506565 352610 506631 352613
rect 248708 352608 506631 352610
rect 248708 352552 506570 352608
rect 506626 352552 506631 352608
rect 248708 352550 506631 352552
rect 248708 352548 248714 352550
rect 506565 352547 506631 352550
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 175273 351114 175339 351117
rect 224166 351114 224172 351116
rect 175273 351112 224172 351114
rect 175273 351056 175278 351112
rect 175334 351056 224172 351112
rect 175273 351054 224172 351056
rect 175273 351051 175339 351054
rect 224166 351052 224172 351054
rect 224236 351052 224242 351116
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2773 306234 2839 306237
rect -960 306232 2839 306234
rect -960 306176 2778 306232
rect 2834 306176 2839 306232
rect -960 306174 2839 306176
rect -960 306084 480 306174
rect 2773 306171 2839 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 202086 254010 202092 254012
rect 6870 253950 202092 254010
rect 202086 253948 202092 253950
rect 202156 253948 202162 254012
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3877 241090 3943 241093
rect -960 241088 3943 241090
rect -960 241032 3882 241088
rect 3938 241032 3943 241088
rect -960 241030 3943 241032
rect -960 240940 480 241030
rect 3877 241027 3943 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3049 214978 3115 214981
rect -960 214976 3115 214978
rect -960 214920 3054 214976
rect 3110 214920 3115 214976
rect -960 214918 3115 214920
rect -960 214828 480 214918
rect 3049 214915 3115 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3785 188866 3851 188869
rect -960 188864 3851 188866
rect -960 188808 3790 188864
rect 3846 188808 3851 188864
rect -960 188806 3851 188808
rect -960 188716 480 188806
rect 3785 188803 3851 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 120073 177714 120139 177717
rect 219750 177714 219756 177716
rect 120073 177712 219756 177714
rect 120073 177656 120078 177712
rect 120134 177656 219756 177712
rect 120073 177654 219756 177656
rect 120073 177651 120139 177654
rect 219750 177652 219756 177654
rect 219820 177652 219826 177716
rect 63493 177578 63559 177581
rect 215518 177578 215524 177580
rect 63493 177576 215524 177578
rect 63493 177520 63498 177576
rect 63554 177520 215524 177576
rect 63493 177518 215524 177520
rect 63493 177515 63559 177518
rect 215518 177516 215524 177518
rect 215588 177516 215594 177580
rect 49693 177442 49759 177445
rect 214414 177442 214420 177444
rect 49693 177440 214420 177442
rect 49693 177384 49698 177440
rect 49754 177384 214420 177440
rect 49693 177382 214420 177384
rect 49693 177379 49759 177382
rect 214414 177380 214420 177382
rect 214484 177380 214490 177444
rect 13813 177306 13879 177309
rect 211470 177306 211476 177308
rect 13813 177304 211476 177306
rect 13813 177248 13818 177304
rect 13874 177248 211476 177304
rect 13813 177246 211476 177248
rect 13813 177243 13879 177246
rect 211470 177244 211476 177246
rect 211540 177244 211546 177308
rect 230606 177244 230612 177308
rect 230676 177306 230682 177308
rect 273253 177306 273319 177309
rect 230676 177304 273319 177306
rect 230676 177248 273258 177304
rect 273314 177248 273319 177304
rect 230676 177246 273319 177248
rect 230676 177244 230682 177246
rect 273253 177243 273319 177246
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3049 162890 3115 162893
rect -960 162888 3115 162890
rect -960 162832 3054 162888
rect 3110 162832 3115 162888
rect -960 162830 3115 162832
rect -960 162740 480 162830
rect 3049 162827 3115 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 254710 87484 254716 87548
rect 254780 87546 254786 87548
rect 576853 87546 576919 87549
rect 254780 87544 576919 87546
rect 254780 87488 576858 87544
rect 576914 87488 576919 87544
rect 254780 87486 576919 87488
rect 254780 87484 254786 87486
rect 576853 87483 576919 87486
rect 234102 86260 234108 86324
rect 234172 86322 234178 86324
rect 307753 86322 307819 86325
rect 234172 86320 307819 86322
rect 234172 86264 307758 86320
rect 307814 86264 307819 86320
rect 234172 86262 307819 86264
rect 234172 86260 234178 86262
rect 307753 86259 307819 86262
rect 248822 86124 248828 86188
rect 248892 86186 248898 86188
rect 503713 86186 503779 86189
rect 248892 86184 503779 86186
rect 248892 86128 503718 86184
rect 503774 86128 503779 86184
rect 248892 86126 503779 86128
rect 248892 86124 248898 86126
rect 503713 86123 503779 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 236862 84764 236868 84828
rect 236932 84826 236938 84828
rect 343633 84826 343699 84829
rect 236932 84824 343699 84826
rect 236932 84768 343638 84824
rect 343694 84768 343699 84824
rect 236932 84766 343699 84768
rect 236932 84764 236938 84766
rect 343633 84763 343699 84766
rect 3601 84690 3667 84693
rect -960 84688 3667 84690
rect -960 84632 3606 84688
rect 3662 84632 3667 84688
rect -960 84630 3667 84632
rect -960 84540 480 84630
rect 3601 84627 3667 84630
rect 241094 82044 241100 82108
rect 241164 82106 241170 82108
rect 398925 82106 398991 82109
rect 241164 82104 398991 82106
rect 241164 82048 398930 82104
rect 398986 82048 398991 82104
rect 241164 82046 398991 82048
rect 241164 82044 241170 82046
rect 398925 82043 398991 82046
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3550 45522 3556 45524
rect -960 45462 3556 45522
rect -960 45372 480 45462
rect 3550 45460 3556 45462
rect 3620 45460 3626 45524
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 264094 31724 264100 31788
rect 264164 31786 264170 31788
rect 583526 31786 583586 32950
rect 264164 31726 583586 31786
rect 264164 31724 264170 31726
rect 247902 26828 247908 26892
rect 247972 26890 247978 26892
rect 487153 26890 487219 26893
rect 247972 26888 487219 26890
rect 247972 26832 487158 26888
rect 487214 26832 487219 26888
rect 247972 26830 487219 26832
rect 247972 26828 247978 26830
rect 487153 26827 487219 26830
rect 235390 25604 235396 25668
rect 235460 25666 235466 25668
rect 325693 25666 325759 25669
rect 235460 25664 325759 25666
rect 235460 25608 325698 25664
rect 325754 25608 325759 25664
rect 235460 25606 325759 25608
rect 235460 25604 235466 25606
rect 325693 25603 325759 25606
rect 254894 25468 254900 25532
rect 254964 25530 254970 25532
rect 574093 25530 574159 25533
rect 254964 25528 574159 25530
rect 254964 25472 574098 25528
rect 574154 25472 574159 25528
rect 254964 25470 574159 25472
rect 254964 25468 254970 25470
rect 574093 25467 574159 25470
rect 243854 24380 243860 24444
rect 243924 24442 243930 24444
rect 432045 24442 432111 24445
rect 243924 24440 432111 24442
rect 243924 24384 432050 24440
rect 432106 24384 432111 24440
rect 243924 24382 432111 24384
rect 243924 24380 243930 24382
rect 432045 24379 432111 24382
rect 246430 24244 246436 24308
rect 246500 24306 246506 24308
rect 466453 24306 466519 24309
rect 246500 24304 466519 24306
rect 246500 24248 466458 24304
rect 466514 24248 466519 24304
rect 246500 24246 466519 24248
rect 246500 24244 246506 24246
rect 466453 24243 466519 24246
rect 246614 24108 246620 24172
rect 246684 24170 246690 24172
rect 470593 24170 470659 24173
rect 246684 24168 470659 24170
rect 246684 24112 470598 24168
rect 470654 24112 470659 24168
rect 246684 24110 470659 24112
rect 246684 24108 246690 24110
rect 470593 24107 470659 24110
rect 239438 22884 239444 22948
rect 239508 22946 239514 22948
rect 382365 22946 382431 22949
rect 239508 22944 382431 22946
rect 239508 22888 382370 22944
rect 382426 22888 382431 22944
rect 239508 22886 382431 22888
rect 239508 22884 239514 22886
rect 382365 22883 382431 22886
rect 242198 22748 242204 22812
rect 242268 22810 242274 22812
rect 414013 22810 414079 22813
rect 242268 22808 414079 22810
rect 242268 22752 414018 22808
rect 414074 22752 414079 22808
rect 242268 22750 414079 22752
rect 242268 22748 242274 22750
rect 414013 22747 414079 22750
rect 242382 22612 242388 22676
rect 242452 22674 242458 22676
rect 416773 22674 416839 22677
rect 242452 22672 416839 22674
rect 242452 22616 416778 22672
rect 416834 22616 416839 22672
rect 242452 22614 416839 22616
rect 242452 22612 242458 22614
rect 416773 22611 416839 22614
rect 237046 21524 237052 21588
rect 237116 21586 237122 21588
rect 346393 21586 346459 21589
rect 237116 21584 346459 21586
rect 237116 21528 346398 21584
rect 346454 21528 346459 21584
rect 237116 21526 346459 21528
rect 237116 21524 237122 21526
rect 346393 21523 346459 21526
rect 238334 21388 238340 21452
rect 238404 21450 238410 21452
rect 360193 21450 360259 21453
rect 238404 21448 360259 21450
rect 238404 21392 360198 21448
rect 360254 21392 360259 21448
rect 238404 21390 360259 21392
rect 238404 21388 238410 21390
rect 360193 21387 360259 21390
rect 239622 21252 239628 21316
rect 239692 21314 239698 21316
rect 378133 21314 378199 21317
rect 239692 21312 378199 21314
rect 239692 21256 378138 21312
rect 378194 21256 378199 21312
rect 239692 21254 378199 21256
rect 239692 21252 239698 21254
rect 378133 21251 378199 21254
rect 232814 20164 232820 20228
rect 232884 20226 232890 20228
rect 289813 20226 289879 20229
rect 232884 20224 289879 20226
rect 232884 20168 289818 20224
rect 289874 20168 289879 20224
rect 232884 20166 289879 20168
rect 232884 20164 232890 20166
rect 289813 20163 289879 20166
rect 232630 20028 232636 20092
rect 232700 20090 232706 20092
rect 292573 20090 292639 20093
rect 232700 20088 292639 20090
rect 232700 20032 292578 20088
rect 292634 20032 292639 20088
rect 232700 20030 292639 20032
rect 232700 20028 232706 20030
rect 292573 20027 292639 20030
rect 234286 19892 234292 19956
rect 234356 19954 234362 19956
rect 307845 19954 307911 19957
rect 234356 19952 307911 19954
rect 234356 19896 307850 19952
rect 307906 19896 307911 19952
rect 234356 19894 307911 19896
rect 234356 19892 234362 19894
rect 307845 19891 307911 19894
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 295926 19348 295932 19412
rect 295996 19410 296002 19412
rect 583526 19410 583586 19622
rect 295996 19350 583586 19410
rect 295996 19348 296002 19350
rect 230790 18532 230796 18596
rect 230860 18594 230866 18596
rect 276105 18594 276171 18597
rect 230860 18592 276171 18594
rect 230860 18536 276110 18592
rect 276166 18536 276171 18592
rect 230860 18534 276171 18536
rect 230860 18532 230866 18534
rect 276105 18531 276171 18534
rect 251950 17444 251956 17508
rect 252020 17506 252026 17508
rect 540973 17506 541039 17509
rect 252020 17504 541039 17506
rect 252020 17448 540978 17504
rect 541034 17448 541039 17504
rect 252020 17446 541039 17448
rect 252020 17444 252026 17446
rect 540973 17443 541039 17446
rect 253238 17308 253244 17372
rect 253308 17370 253314 17372
rect 556245 17370 556311 17373
rect 253308 17368 556311 17370
rect 253308 17312 556250 17368
rect 556306 17312 556311 17368
rect 253308 17310 556311 17312
rect 253308 17308 253314 17310
rect 556245 17307 556311 17310
rect 253422 17172 253428 17236
rect 253492 17234 253498 17236
rect 558913 17234 558979 17237
rect 253492 17232 558979 17234
rect 253492 17176 558918 17232
rect 558974 17176 558979 17232
rect 253492 17174 558979 17176
rect 253492 17172 253498 17174
rect 558913 17171 558979 17174
rect 138841 16010 138907 16013
rect 221038 16010 221044 16012
rect 138841 16008 221044 16010
rect 138841 15952 138846 16008
rect 138902 15952 221044 16008
rect 138841 15950 221044 15952
rect 138841 15947 138907 15950
rect 221038 15948 221044 15950
rect 221108 15948 221114 16012
rect 250846 15948 250852 16012
rect 250916 16010 250922 16012
rect 520273 16010 520339 16013
rect 250916 16008 520339 16010
rect 250916 15952 520278 16008
rect 520334 15952 520339 16008
rect 250916 15950 520339 15952
rect 250916 15948 250922 15950
rect 520273 15947 520339 15950
rect 84193 15874 84259 15877
rect 217174 15874 217180 15876
rect 84193 15872 217180 15874
rect 84193 15816 84198 15872
rect 84254 15816 217180 15872
rect 84193 15814 217180 15816
rect 84193 15811 84259 15814
rect 217174 15812 217180 15814
rect 217244 15812 217250 15876
rect 250662 15812 250668 15876
rect 250732 15874 250738 15876
rect 523769 15874 523835 15877
rect 250732 15872 523835 15874
rect 250732 15816 523774 15872
rect 523830 15816 523835 15872
rect 250732 15814 523835 15816
rect 250732 15812 250738 15814
rect 523769 15811 523835 15814
rect 155217 14786 155283 14789
rect 218830 14786 218836 14788
rect 155217 14784 218836 14786
rect 155217 14728 155222 14784
rect 155278 14728 218836 14784
rect 155217 14726 218836 14728
rect 155217 14723 155283 14726
rect 218830 14724 218836 14726
rect 218900 14724 218906 14788
rect 246798 14724 246804 14788
rect 246868 14786 246874 14788
rect 469857 14786 469923 14789
rect 246868 14784 469923 14786
rect 246868 14728 469862 14784
rect 469918 14728 469923 14784
rect 246868 14726 469923 14728
rect 246868 14724 246874 14726
rect 469857 14723 469923 14726
rect 81617 14650 81683 14653
rect 216990 14650 216996 14652
rect 81617 14648 216996 14650
rect 81617 14592 81622 14648
rect 81678 14592 216996 14648
rect 81617 14590 216996 14592
rect 81617 14587 81683 14590
rect 216990 14588 216996 14590
rect 217060 14588 217066 14652
rect 248270 14588 248276 14652
rect 248340 14650 248346 14652
rect 484761 14650 484827 14653
rect 248340 14648 484827 14650
rect 248340 14592 484766 14648
rect 484822 14592 484827 14648
rect 248340 14590 484827 14592
rect 248340 14588 248346 14590
rect 484761 14587 484827 14590
rect 13537 14514 13603 14517
rect 211286 14514 211292 14516
rect 13537 14512 211292 14514
rect 13537 14456 13542 14512
rect 13598 14456 211292 14512
rect 13537 14454 211292 14456
rect 13537 14451 13603 14454
rect 211286 14452 211292 14454
rect 211356 14452 211362 14516
rect 248086 14452 248092 14516
rect 248156 14514 248162 14516
rect 488809 14514 488875 14517
rect 248156 14512 488875 14514
rect 248156 14456 488814 14512
rect 488870 14456 488875 14512
rect 248156 14454 488875 14456
rect 248156 14452 248162 14454
rect 488809 14451 488875 14454
rect 66713 13154 66779 13157
rect 215702 13154 215708 13156
rect 66713 13152 215708 13154
rect 66713 13096 66718 13152
rect 66774 13096 215708 13152
rect 66713 13094 215708 13096
rect 66713 13091 66779 13094
rect 215702 13092 215708 13094
rect 215772 13092 215778 13156
rect 244038 13092 244044 13156
rect 244108 13154 244114 13156
rect 433977 13154 434043 13157
rect 244108 13152 434043 13154
rect 244108 13096 433982 13152
rect 434038 13096 434043 13152
rect 244108 13094 434043 13096
rect 244108 13092 244114 13094
rect 433977 13091 434043 13094
rect 48497 13018 48563 13021
rect 214230 13018 214236 13020
rect 48497 13016 214236 13018
rect 48497 12960 48502 13016
rect 48558 12960 214236 13016
rect 48497 12958 214236 12960
rect 48497 12955 48563 12958
rect 214230 12956 214236 12958
rect 214300 12956 214306 13020
rect 245510 12956 245516 13020
rect 245580 13018 245586 13020
rect 451641 13018 451707 13021
rect 245580 13016 451707 13018
rect 245580 12960 451646 13016
rect 451702 12960 451707 13016
rect 245580 12958 451707 12960
rect 245580 12956 245586 12958
rect 451641 12955 451707 12958
rect 122281 11930 122347 11933
rect 219566 11930 219572 11932
rect 122281 11928 219572 11930
rect 122281 11872 122286 11928
rect 122342 11872 219572 11928
rect 122281 11870 219572 11872
rect 122281 11867 122347 11870
rect 219566 11868 219572 11870
rect 219636 11868 219642 11932
rect 118785 11794 118851 11797
rect 219198 11794 219204 11796
rect 118785 11792 219204 11794
rect 118785 11736 118790 11792
rect 118846 11736 219204 11792
rect 118785 11734 219204 11736
rect 118785 11731 118851 11734
rect 219198 11732 219204 11734
rect 219268 11732 219274 11796
rect 242750 11732 242756 11796
rect 242820 11794 242826 11796
rect 412633 11794 412699 11797
rect 242820 11792 412699 11794
rect 242820 11736 412638 11792
rect 412694 11736 412699 11792
rect 242820 11734 412699 11736
rect 242820 11732 242826 11734
rect 412633 11731 412699 11734
rect 17033 11658 17099 11661
rect 211102 11658 211108 11660
rect 17033 11656 211108 11658
rect 17033 11600 17038 11656
rect 17094 11600 211108 11656
rect 17033 11598 211108 11600
rect 17033 11595 17099 11598
rect 211102 11596 211108 11598
rect 211172 11596 211178 11660
rect 242566 11596 242572 11660
rect 242636 11658 242642 11660
rect 415485 11658 415551 11661
rect 242636 11656 415551 11658
rect 242636 11600 415490 11656
rect 415546 11600 415551 11656
rect 242636 11598 415551 11600
rect 242636 11596 242642 11598
rect 415485 11595 415551 11598
rect 100753 10570 100819 10573
rect 218646 10570 218652 10572
rect 100753 10568 218652 10570
rect 100753 10512 100758 10568
rect 100814 10512 218652 10568
rect 100753 10510 218652 10512
rect 100753 10507 100819 10510
rect 218646 10508 218652 10510
rect 218716 10508 218722 10572
rect 237966 10508 237972 10572
rect 238036 10570 238042 10572
rect 363505 10570 363571 10573
rect 238036 10568 363571 10570
rect 238036 10512 363510 10568
rect 363566 10512 363571 10568
rect 238036 10510 363571 10512
rect 238036 10508 238042 10510
rect 363505 10507 363571 10510
rect 86401 10434 86467 10437
rect 216622 10434 216628 10436
rect 86401 10432 216628 10434
rect 86401 10376 86406 10432
rect 86462 10376 216628 10432
rect 86401 10374 216628 10376
rect 86401 10371 86467 10374
rect 216622 10372 216628 10374
rect 216692 10372 216698 10436
rect 239806 10372 239812 10436
rect 239876 10434 239882 10436
rect 377673 10434 377739 10437
rect 239876 10432 377739 10434
rect 239876 10376 377678 10432
rect 377734 10376 377739 10432
rect 239876 10374 377739 10376
rect 239876 10372 239882 10374
rect 377673 10371 377739 10374
rect 83273 10298 83339 10301
rect 216806 10298 216812 10300
rect 83273 10296 216812 10298
rect 83273 10240 83278 10296
rect 83334 10240 216812 10296
rect 83273 10238 216812 10240
rect 83273 10235 83339 10238
rect 216806 10236 216812 10238
rect 216876 10236 216882 10300
rect 239990 10236 239996 10300
rect 240060 10298 240066 10300
rect 381169 10298 381235 10301
rect 240060 10296 381235 10298
rect 240060 10240 381174 10296
rect 381230 10240 381235 10296
rect 240060 10238 381235 10240
rect 240060 10236 240066 10238
rect 381169 10235 381235 10238
rect 235574 9148 235580 9212
rect 235644 9210 235650 9212
rect 327993 9210 328059 9213
rect 235644 9208 328059 9210
rect 235644 9152 327998 9208
rect 328054 9152 328059 9208
rect 235644 9150 328059 9152
rect 235644 9148 235650 9150
rect 327993 9147 328059 9150
rect 51349 9074 51415 9077
rect 214046 9074 214052 9076
rect 51349 9072 214052 9074
rect 51349 9016 51354 9072
rect 51410 9016 214052 9072
rect 51349 9014 214052 9016
rect 51349 9011 51415 9014
rect 214046 9012 214052 9014
rect 214116 9012 214122 9076
rect 237230 9012 237236 9076
rect 237300 9074 237306 9076
rect 345749 9074 345815 9077
rect 237300 9072 345815 9074
rect 237300 9016 345754 9072
rect 345810 9016 345815 9072
rect 237300 9014 345815 9016
rect 237300 9012 237306 9014
rect 345749 9011 345815 9014
rect 565 8938 631 8941
rect 209814 8938 209820 8940
rect 565 8936 209820 8938
rect 565 8880 570 8936
rect 626 8880 209820 8936
rect 565 8878 209820 8880
rect 565 8875 631 8878
rect 209814 8876 209820 8878
rect 209884 8876 209890 8940
rect 252134 8876 252140 8940
rect 252204 8938 252210 8940
rect 539593 8938 539659 8941
rect 252204 8936 539659 8938
rect 252204 8880 539598 8936
rect 539654 8880 539659 8936
rect 252204 8878 539659 8880
rect 252204 8876 252210 8878
rect 539593 8875 539659 8878
rect 206185 7986 206251 7989
rect 226374 7986 226380 7988
rect 206185 7984 226380 7986
rect 206185 7928 206190 7984
rect 206246 7928 226380 7984
rect 206185 7926 226380 7928
rect 206185 7923 206251 7926
rect 226374 7924 226380 7926
rect 226444 7924 226450 7988
rect 192017 7850 192083 7853
rect 225270 7850 225276 7852
rect 192017 7848 225276 7850
rect 192017 7792 192022 7848
rect 192078 7792 225276 7848
rect 192017 7790 225276 7792
rect 192017 7787 192083 7790
rect 225270 7788 225276 7790
rect 225340 7788 225346 7852
rect 174261 7714 174327 7717
rect 223982 7714 223988 7716
rect 174261 7712 223988 7714
rect 174261 7656 174266 7712
rect 174322 7656 223988 7712
rect 174261 7654 223988 7656
rect 174261 7651 174327 7654
rect 223982 7652 223988 7654
rect 224052 7652 224058 7716
rect 170765 7578 170831 7581
rect 223798 7578 223804 7580
rect 170765 7576 223804 7578
rect 170765 7520 170770 7576
rect 170826 7520 223804 7576
rect 170765 7518 223804 7520
rect 170765 7515 170831 7518
rect 223798 7516 223804 7518
rect 223868 7516 223874 7580
rect 233918 7516 233924 7580
rect 233988 7578 233994 7580
rect 310237 7578 310303 7581
rect 233988 7576 310303 7578
rect 233988 7520 310242 7576
rect 310298 7520 310303 7576
rect 233988 7518 310303 7520
rect 233988 7516 233994 7518
rect 310237 7515 310303 7518
rect 194409 6626 194475 6629
rect 224902 6626 224908 6628
rect 194409 6624 224908 6626
rect -960 6490 480 6580
rect 194409 6568 194414 6624
rect 194470 6568 224908 6624
rect 194409 6566 224908 6568
rect 194409 6563 194475 6566
rect 224902 6564 224908 6566
rect 224972 6564 224978 6628
rect 583520 6626 584960 6716
rect 583342 6566 584960 6626
rect 3366 6490 3372 6492
rect -960 6430 3372 6490
rect -960 6340 480 6430
rect 3366 6428 3372 6430
rect 3436 6428 3442 6492
rect 190821 6490 190887 6493
rect 225086 6490 225092 6492
rect 190821 6488 225092 6490
rect 190821 6432 190826 6488
rect 190882 6432 225092 6488
rect 190821 6430 225092 6432
rect 190821 6427 190887 6430
rect 225086 6428 225092 6430
rect 225156 6428 225162 6492
rect 230974 6428 230980 6492
rect 231044 6490 231050 6492
rect 274817 6490 274883 6493
rect 231044 6488 274883 6490
rect 231044 6432 274822 6488
rect 274878 6432 274883 6488
rect 231044 6430 274883 6432
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect 231044 6428 231050 6430
rect 274817 6427 274883 6430
rect 173157 6354 173223 6357
rect 223614 6354 223620 6356
rect 173157 6352 223620 6354
rect 173157 6296 173162 6352
rect 173218 6296 223620 6352
rect 173157 6294 223620 6296
rect 173157 6291 173223 6294
rect 223614 6292 223620 6294
rect 223684 6292 223690 6356
rect 232998 6292 233004 6356
rect 233068 6354 233074 6356
rect 292573 6354 292639 6357
rect 233068 6352 292639 6354
rect 233068 6296 292578 6352
rect 292634 6296 292639 6352
rect 233068 6294 292639 6296
rect 233068 6292 233074 6294
rect 292573 6291 292639 6294
rect 137645 6218 137711 6221
rect 220854 6218 220860 6220
rect 137645 6216 220860 6218
rect 137645 6160 137650 6216
rect 137706 6160 220860 6216
rect 137645 6158 220860 6160
rect 137645 6155 137711 6158
rect 220854 6156 220860 6158
rect 220924 6156 220930 6220
rect 255078 6156 255084 6220
rect 255148 6218 255154 6220
rect 576301 6218 576367 6221
rect 255148 6216 576367 6218
rect 255148 6160 576306 6216
rect 576362 6160 576367 6216
rect 255148 6158 576367 6160
rect 255148 6156 255154 6158
rect 576301 6155 576367 6158
rect 298502 5612 298508 5676
rect 298572 5674 298578 5676
rect 583526 5674 583586 6430
rect 298572 5614 583586 5674
rect 298572 5612 298578 5614
rect 229870 5340 229876 5404
rect 229940 5402 229946 5404
rect 237373 5402 237439 5405
rect 229940 5400 237439 5402
rect 229940 5344 237378 5400
rect 237434 5344 237439 5400
rect 229940 5342 237439 5344
rect 229940 5340 229946 5342
rect 237373 5339 237439 5342
rect 230054 5204 230060 5268
rect 230124 5266 230130 5268
rect 254669 5266 254735 5269
rect 230124 5264 254735 5266
rect 230124 5208 254674 5264
rect 254730 5208 254735 5264
rect 230124 5206 254735 5208
rect 230124 5204 230130 5206
rect 254669 5203 254735 5206
rect 251030 5068 251036 5132
rect 251100 5130 251106 5132
rect 523033 5130 523099 5133
rect 251100 5128 523099 5130
rect 251100 5072 523038 5128
rect 523094 5072 523099 5128
rect 251100 5070 523099 5072
rect 251100 5068 251106 5070
rect 523033 5067 523099 5070
rect 252318 4932 252324 4996
rect 252388 4994 252394 4996
rect 540789 4994 540855 4997
rect 252388 4992 540855 4994
rect 252388 4936 540794 4992
rect 540850 4936 540855 4992
rect 252388 4934 540855 4936
rect 252388 4932 252394 4934
rect 540789 4931 540855 4934
rect 253606 4796 253612 4860
rect 253676 4858 253682 4860
rect 558545 4858 558611 4861
rect 253676 4856 558611 4858
rect 253676 4800 558550 4856
rect 558606 4800 558611 4856
rect 253676 4798 558611 4800
rect 253676 4796 253682 4798
rect 558545 4795 558611 4798
rect 228950 3708 228956 3772
rect 229020 3770 229026 3772
rect 239305 3770 239371 3773
rect 229020 3768 239371 3770
rect 229020 3712 239310 3768
rect 239366 3712 239371 3768
rect 229020 3710 239371 3712
rect 229020 3708 229026 3710
rect 239305 3707 239371 3710
rect 228582 3572 228588 3636
rect 228652 3634 228658 3636
rect 240501 3634 240567 3637
rect 228652 3632 240567 3634
rect 228652 3576 240506 3632
rect 240562 3576 240567 3632
rect 228652 3574 240567 3576
rect 228652 3572 228658 3574
rect 240501 3571 240567 3574
rect 228766 3436 228772 3500
rect 228836 3498 228842 3500
rect 242893 3498 242959 3501
rect 228836 3496 242959 3498
rect 228836 3440 242898 3496
rect 242954 3440 242959 3496
rect 228836 3438 242959 3440
rect 228836 3436 228842 3438
rect 242893 3435 242959 3438
rect 249006 3436 249012 3500
rect 249076 3498 249082 3500
rect 505369 3498 505435 3501
rect 249076 3496 505435 3498
rect 249076 3440 505374 3496
rect 505430 3440 505435 3496
rect 249076 3438 505435 3440
rect 249076 3436 249082 3438
rect 505369 3435 505435 3438
rect 230238 3300 230244 3364
rect 230308 3362 230314 3364
rect 257061 3362 257127 3365
rect 230308 3360 257127 3362
rect 230308 3304 257066 3360
rect 257122 3304 257127 3360
rect 230308 3302 257127 3304
rect 230308 3300 230314 3302
rect 257061 3299 257127 3302
rect 262622 3300 262628 3364
rect 262692 3362 262698 3364
rect 579797 3362 579863 3365
rect 262692 3360 579863 3362
rect 262692 3304 579802 3360
rect 579858 3304 579863 3360
rect 262692 3302 579863 3304
rect 262692 3300 262698 3302
rect 579797 3299 579863 3302
<< via3 >>
rect 102364 597484 102428 597548
rect 105308 597484 105372 597548
rect 207612 597484 207676 597548
rect 208900 597484 208964 597548
rect 210004 597544 210068 597548
rect 210004 597488 210054 597544
rect 210054 597488 210068 597544
rect 210004 597484 210068 597488
rect 211108 597544 211172 597548
rect 211108 597488 211158 597544
rect 211158 597488 211172 597544
rect 211108 597484 211172 597488
rect 212396 597544 212460 597548
rect 212396 597488 212446 597544
rect 212446 597488 212460 597544
rect 212396 597484 212460 597488
rect 213500 597484 213564 597548
rect 214788 597544 214852 597548
rect 214788 597488 214838 597544
rect 214838 597488 214852 597544
rect 214788 597484 214852 597488
rect 215340 597544 215404 597548
rect 215340 597488 215354 597544
rect 215354 597488 215404 597544
rect 215340 597484 215404 597488
rect 215708 597484 215772 597548
rect 225460 597484 225524 597548
rect 235580 597484 235644 597548
rect 245516 597544 245580 597548
rect 245516 597488 245566 597544
rect 245566 597488 245580 597544
rect 245516 597484 245580 597488
rect 250484 597484 250548 597548
rect 317644 597484 317708 597548
rect 318932 597484 318996 597548
rect 320036 597544 320100 597548
rect 320036 597488 320086 597544
rect 320086 597488 320100 597544
rect 320036 597484 320100 597488
rect 321140 597484 321204 597548
rect 322244 597544 322308 597548
rect 322244 597488 322294 597544
rect 322294 597488 322308 597544
rect 322244 597484 322308 597488
rect 323348 597484 323412 597548
rect 325188 597484 325252 597548
rect 325740 597544 325804 597548
rect 325740 597488 325790 597544
rect 325790 597488 325804 597544
rect 325740 597484 325804 597488
rect 330524 597484 330588 597548
rect 345612 597484 345676 597548
rect 360516 597484 360580 597548
rect 440372 597484 440436 597548
rect 450492 597484 450556 597548
rect 460428 597484 460492 597548
rect 92980 597348 93044 597412
rect 98868 597348 98932 597412
rect 101076 597348 101140 597412
rect 324820 597348 324884 597412
rect 435588 597348 435652 597412
rect 103284 597212 103348 597276
rect 105676 597212 105740 597276
rect 230612 597212 230676 597276
rect 422892 597212 422956 597276
rect 427676 597212 427740 597276
rect 428964 597212 429028 597276
rect 430988 597212 431052 597276
rect 99972 597076 100036 597140
rect 104756 597136 104820 597140
rect 104756 597080 104806 597136
rect 104806 597080 104820 597136
rect 104756 597076 104820 597080
rect 205404 597076 205468 597140
rect 350396 597076 350460 597140
rect 429884 597076 429948 597140
rect 94268 596940 94332 597004
rect 97764 596940 97828 597004
rect 130516 596940 130580 597004
rect 315252 596940 315316 597004
rect 340460 596940 340524 597004
rect 424180 596940 424244 597004
rect 431724 596940 431788 597004
rect 433380 597000 433444 597004
rect 433380 596944 433394 597000
rect 433394 596944 433444 597000
rect 433380 596940 433444 596944
rect 434668 597000 434732 597004
rect 434668 596944 434718 597000
rect 434718 596944 434732 597000
rect 434668 596940 434732 596944
rect 110460 596804 110524 596868
rect 240548 596804 240612 596868
rect 314332 596804 314396 596868
rect 465396 596804 465460 596868
rect 125548 596668 125612 596732
rect 435220 596668 435284 596732
rect 445524 596668 445588 596732
rect 135484 596532 135548 596596
rect 140636 596592 140700 596596
rect 140636 596536 140686 596592
rect 140686 596536 140700 596592
rect 140636 596532 140700 596536
rect 312860 596532 312924 596596
rect 202828 596456 202892 596460
rect 202828 596400 202878 596456
rect 202878 596400 202892 596456
rect 202828 596396 202892 596400
rect 425284 596396 425348 596460
rect 95372 596260 95436 596324
rect 115612 596260 115676 596324
rect 120580 596260 120644 596324
rect 204300 596320 204364 596324
rect 204300 596264 204314 596320
rect 204314 596264 204364 596320
rect 204300 596260 204364 596264
rect 219204 596260 219268 596324
rect 335124 596260 335188 596324
rect 354444 596260 354508 596324
rect 455460 596320 455524 596324
rect 455460 596264 455474 596320
rect 455474 596264 455524 596320
rect 455460 596260 455524 596264
rect 470364 596260 470428 596324
rect 282132 589868 282196 589932
rect 407804 526628 407868 526692
rect 407620 523636 407684 523700
rect 407620 489772 407684 489836
rect 92980 488472 93044 488476
rect 92980 488416 92994 488472
rect 92994 488416 93044 488472
rect 92980 488412 93044 488416
rect 94268 488472 94332 488476
rect 94268 488416 94282 488472
rect 94282 488416 94332 488472
rect 94268 488412 94332 488416
rect 95372 488472 95436 488476
rect 95372 488416 95386 488472
rect 95386 488416 95436 488472
rect 95372 488412 95436 488416
rect 97764 488472 97828 488476
rect 97764 488416 97814 488472
rect 97814 488416 97828 488472
rect 97764 488412 97828 488416
rect 98868 488472 98932 488476
rect 98868 488416 98918 488472
rect 98918 488416 98932 488472
rect 98868 488412 98932 488416
rect 99972 488472 100036 488476
rect 99972 488416 100022 488472
rect 100022 488416 100036 488472
rect 99972 488412 100036 488416
rect 101076 488472 101140 488476
rect 101076 488416 101126 488472
rect 101126 488416 101140 488472
rect 101076 488412 101140 488416
rect 102364 488472 102428 488476
rect 102364 488416 102414 488472
rect 102414 488416 102428 488472
rect 102364 488412 102428 488416
rect 104756 488472 104820 488476
rect 104756 488416 104806 488472
rect 104806 488416 104820 488472
rect 104756 488412 104820 488416
rect 105676 488472 105740 488476
rect 105676 488416 105726 488472
rect 105726 488416 105740 488472
rect 105676 488412 105740 488416
rect 204300 488412 204364 488476
rect 214788 488472 214852 488476
rect 214788 488416 214838 488472
rect 214838 488416 214852 488472
rect 214788 488412 214852 488416
rect 314332 488472 314396 488476
rect 314332 488416 314346 488472
rect 314346 488416 314396 488472
rect 314332 488412 314396 488416
rect 315436 488472 315500 488476
rect 315436 488416 315450 488472
rect 315450 488416 315500 488472
rect 315436 488412 315500 488416
rect 323348 488412 323412 488476
rect 422892 488412 422956 488476
rect 424180 488412 424244 488476
rect 425284 488412 425348 488476
rect 211108 488336 211172 488340
rect 211108 488280 211158 488336
rect 211158 488280 211172 488336
rect 211108 488276 211172 488280
rect 213500 488276 213564 488340
rect 215708 488276 215772 488340
rect 465396 488276 465460 488340
rect 105308 488140 105372 488204
rect 110460 488140 110524 488204
rect 203012 488140 203076 488204
rect 429884 488140 429948 488204
rect 103284 488004 103348 488068
rect 407804 488004 407868 488068
rect 313044 487928 313108 487932
rect 313044 487872 313058 487928
rect 313058 487872 313108 487928
rect 313044 487868 313108 487872
rect 428964 487732 429028 487796
rect 427676 487596 427740 487660
rect 435588 487596 435652 487660
rect 212212 487460 212276 487524
rect 321140 487460 321204 487524
rect 324820 487460 324884 487524
rect 430988 487460 431052 487524
rect 432276 487460 432340 487524
rect 433380 487520 433444 487524
rect 433380 487464 433394 487520
rect 433394 487464 433444 487520
rect 433380 487460 433444 487464
rect 434852 487460 434916 487524
rect 210004 487324 210068 487388
rect 318932 487324 318996 487388
rect 115612 487188 115676 487252
rect 120580 487188 120644 487252
rect 125548 487188 125612 487252
rect 130516 487188 130580 487252
rect 135484 487188 135548 487252
rect 140636 487248 140700 487252
rect 140636 487192 140686 487248
rect 140686 487192 140700 487248
rect 140636 487188 140700 487192
rect 203012 487188 203076 487252
rect 205404 487188 205468 487252
rect 207612 487248 207676 487252
rect 207612 487192 207662 487248
rect 207662 487192 207676 487248
rect 207612 487188 207676 487192
rect 208900 487188 208964 487252
rect 215340 487188 215404 487252
rect 220492 487188 220556 487252
rect 225460 487188 225524 487252
rect 230612 487188 230676 487252
rect 235580 487188 235644 487252
rect 240548 487188 240612 487252
rect 245516 487188 245580 487252
rect 250484 487188 250548 487252
rect 317644 487188 317708 487252
rect 320036 487248 320100 487252
rect 320036 487192 320086 487248
rect 320086 487192 320100 487248
rect 320036 487188 320100 487192
rect 322244 487248 322308 487252
rect 322244 487192 322258 487248
rect 322258 487192 322308 487248
rect 322244 487188 322308 487192
rect 325188 487188 325252 487252
rect 325740 487188 325804 487252
rect 330524 487188 330588 487252
rect 335492 487188 335556 487252
rect 340460 487188 340524 487252
rect 345612 487188 345676 487252
rect 350396 487188 350460 487252
rect 355548 487188 355612 487252
rect 360516 487188 360580 487252
rect 435220 487188 435284 487252
rect 440372 487188 440436 487252
rect 445524 487188 445588 487252
rect 450492 487188 450556 487252
rect 455460 487188 455524 487252
rect 460428 487188 460492 487252
rect 470732 487188 470796 487252
rect 382228 454276 382292 454340
rect 378732 454140 378796 454204
rect 379100 454004 379164 454068
rect 3556 446796 3620 446860
rect 202092 446524 202156 446588
rect 3372 446388 3436 446452
rect 282132 446388 282196 446452
rect 298508 446388 298572 446452
rect 264284 445844 264348 445908
rect 262628 445708 262692 445772
rect 262812 445028 262876 445092
rect 295932 444348 295996 444412
rect 211844 444076 211908 444140
rect 212396 444076 212460 444140
rect 212948 444076 213012 444140
rect 251036 444076 251100 444140
rect 256556 444076 256620 444140
rect 264100 443532 264164 443596
rect 251036 442716 251100 442780
rect 256556 442580 256620 442644
rect 212948 442444 213012 442508
rect 211844 442308 211908 442372
rect 212396 442172 212460 442236
rect 383332 425716 383396 425780
rect 332548 400964 332612 401028
rect 332548 400616 332612 400620
rect 332548 400560 332598 400616
rect 332598 400560 332612 400616
rect 332548 400556 332612 400560
rect 253060 399196 253124 399260
rect 228772 398108 228836 398172
rect 254532 398788 254596 398852
rect 264284 398788 264348 398852
rect 262812 398652 262876 398716
rect 216628 397836 216692 397900
rect 225460 397836 225524 397900
rect 230428 397836 230492 397900
rect 233188 397836 233252 397900
rect 242388 397836 242452 397900
rect 246988 397836 247052 397900
rect 247724 397836 247788 397900
rect 251956 397836 252020 397900
rect 254532 397836 254596 397900
rect 211108 397700 211172 397764
rect 212764 397700 212828 397764
rect 214420 397700 214484 397764
rect 215340 397700 215404 397764
rect 217180 397700 217244 397764
rect 219020 397700 219084 397764
rect 221228 397700 221292 397764
rect 222148 397760 222212 397764
rect 222148 397704 222198 397760
rect 222198 397704 222212 397760
rect 222148 397700 222212 397704
rect 223804 397700 223868 397764
rect 224908 397700 224972 397764
rect 229876 397700 229940 397764
rect 230612 397700 230676 397764
rect 232636 397700 232700 397764
rect 233924 397700 233988 397764
rect 235212 397700 235276 397764
rect 236868 397700 236932 397764
rect 237972 397700 238036 397764
rect 239444 397700 239508 397764
rect 242204 397700 242268 397764
rect 243676 397700 243740 397764
rect 246620 397700 246684 397764
rect 247908 397700 247972 397764
rect 248644 397700 248708 397764
rect 250668 397700 250732 397764
rect 251772 397700 251836 397764
rect 253428 397700 253492 397764
rect 254716 397700 254780 397764
rect 211476 397624 211540 397628
rect 211476 397568 211490 397624
rect 211490 397568 211540 397624
rect 211476 397564 211540 397568
rect 214052 397564 214116 397628
rect 215708 397564 215772 397628
rect 216996 397564 217060 397628
rect 218836 397564 218900 397628
rect 219572 397564 219636 397628
rect 220860 397564 220924 397628
rect 221412 397564 221476 397628
rect 223988 397564 224052 397628
rect 225092 397624 225156 397628
rect 225092 397568 225142 397624
rect 225142 397568 225156 397624
rect 225092 397564 225156 397568
rect 226564 397624 226628 397628
rect 226564 397568 226578 397624
rect 226578 397568 226628 397624
rect 226564 397564 226628 397568
rect 228588 397564 228652 397628
rect 230060 397624 230124 397628
rect 230060 397568 230110 397624
rect 230110 397568 230124 397624
rect 230060 397564 230124 397568
rect 230796 397564 230860 397628
rect 232820 397624 232884 397628
rect 232820 397568 232870 397624
rect 232870 397568 232884 397624
rect 232820 397564 232884 397568
rect 234108 397564 234172 397628
rect 235396 397564 235460 397628
rect 237052 397564 237116 397628
rect 238156 397564 238220 397628
rect 239628 397564 239692 397628
rect 242756 397564 242820 397628
rect 243860 397564 243924 397628
rect 246436 397564 246500 397628
rect 248092 397564 248156 397628
rect 248828 397564 248892 397628
rect 250852 397624 250916 397628
rect 250852 397568 250866 397624
rect 250866 397568 250916 397624
rect 250852 397564 250916 397568
rect 252140 397564 252204 397628
rect 253244 397564 253308 397628
rect 254900 397564 254964 397628
rect 209820 397428 209884 397492
rect 211292 397488 211356 397492
rect 211292 397432 211342 397488
rect 211342 397432 211356 397488
rect 211292 397428 211356 397432
rect 212580 397488 212644 397492
rect 212580 397432 212630 397488
rect 212630 397432 212644 397488
rect 212580 397428 212644 397432
rect 214236 397428 214300 397492
rect 215524 397428 215588 397492
rect 216812 397488 216876 397492
rect 216812 397432 216826 397488
rect 216826 397432 216876 397488
rect 216812 397428 216876 397432
rect 218652 397428 218716 397492
rect 219388 397428 219452 397492
rect 219756 397488 219820 397492
rect 219756 397432 219770 397488
rect 219770 397432 219820 397488
rect 219756 397428 219820 397432
rect 221044 397488 221108 397492
rect 221044 397432 221094 397488
rect 221094 397432 221108 397488
rect 221044 397428 221108 397432
rect 223068 397428 223132 397492
rect 223620 397428 223684 397492
rect 224172 397428 224236 397492
rect 225276 397488 225340 397492
rect 225276 397432 225290 397488
rect 225290 397432 225340 397488
rect 225276 397428 225340 397432
rect 226380 397488 226444 397492
rect 226380 397432 226394 397488
rect 226394 397432 226444 397488
rect 226380 397428 226444 397432
rect 228956 397488 229020 397492
rect 228956 397432 228970 397488
rect 228970 397432 229020 397488
rect 228956 397428 229020 397432
rect 230244 397488 230308 397492
rect 230244 397432 230294 397488
rect 230294 397432 230308 397488
rect 230244 397428 230308 397432
rect 230980 397428 231044 397492
rect 233004 397488 233068 397492
rect 233004 397432 233054 397488
rect 233054 397432 233068 397488
rect 233004 397428 233068 397432
rect 234292 397488 234356 397492
rect 234292 397432 234306 397488
rect 234306 397432 234356 397488
rect 234292 397428 234356 397432
rect 235580 397428 235644 397492
rect 237236 397488 237300 397492
rect 237236 397432 237250 397488
rect 237250 397432 237300 397488
rect 237236 397428 237300 397432
rect 238340 397488 238404 397492
rect 238340 397432 238390 397488
rect 238390 397432 238404 397488
rect 238340 397428 238404 397432
rect 239812 397428 239876 397492
rect 239996 397488 240060 397492
rect 239996 397432 240010 397488
rect 240010 397432 240060 397488
rect 239996 397428 240060 397432
rect 241100 397428 241164 397492
rect 242572 397428 242636 397492
rect 244044 397488 244108 397492
rect 244044 397432 244094 397488
rect 244094 397432 244108 397488
rect 244044 397428 244108 397432
rect 245516 397488 245580 397492
rect 245516 397432 245530 397488
rect 245530 397432 245580 397488
rect 245516 397428 245580 397432
rect 246804 397488 246868 397492
rect 246804 397432 246854 397488
rect 246854 397432 246868 397488
rect 246804 397428 246868 397432
rect 248276 397428 248340 397492
rect 249012 397428 249076 397492
rect 251036 397488 251100 397492
rect 251036 397432 251050 397488
rect 251050 397432 251100 397488
rect 251036 397428 251100 397432
rect 252324 397488 252388 397492
rect 252324 397432 252374 397488
rect 252374 397432 252388 397488
rect 252324 397428 252388 397432
rect 253612 397428 253676 397492
rect 255084 397488 255148 397492
rect 255084 397432 255134 397488
rect 255134 397432 255148 397488
rect 255084 397428 255148 397432
rect 222148 396884 222212 396948
rect 215340 395524 215404 395588
rect 246988 395524 247052 395588
rect 230428 395388 230492 395452
rect 212764 395252 212828 395316
rect 253060 395252 253124 395316
rect 221228 394708 221292 394772
rect 221412 393892 221476 393956
rect 233188 393892 233252 393956
rect 226564 392804 226628 392868
rect 225460 392668 225524 392732
rect 212580 392532 212644 392596
rect 219020 355268 219084 355332
rect 235212 355268 235276 355332
rect 238156 354044 238220 354108
rect 251772 353908 251836 353972
rect 243676 352820 243740 352884
rect 247724 352684 247788 352748
rect 223068 352548 223132 352612
rect 248644 352548 248708 352612
rect 224172 351052 224236 351116
rect 202092 253948 202156 254012
rect 219756 177652 219820 177716
rect 215524 177516 215588 177580
rect 214420 177380 214484 177444
rect 211476 177244 211540 177308
rect 230612 177244 230676 177308
rect 254716 87484 254780 87548
rect 234108 86260 234172 86324
rect 248828 86124 248892 86188
rect 236868 84764 236932 84828
rect 241100 82044 241164 82108
rect 3556 45460 3620 45524
rect 264100 31724 264164 31788
rect 247908 26828 247972 26892
rect 235396 25604 235460 25668
rect 254900 25468 254964 25532
rect 243860 24380 243924 24444
rect 246436 24244 246500 24308
rect 246620 24108 246684 24172
rect 239444 22884 239508 22948
rect 242204 22748 242268 22812
rect 242388 22612 242452 22676
rect 237052 21524 237116 21588
rect 238340 21388 238404 21452
rect 239628 21252 239692 21316
rect 232820 20164 232884 20228
rect 232636 20028 232700 20092
rect 234292 19892 234356 19956
rect 295932 19348 295996 19412
rect 230796 18532 230860 18596
rect 251956 17444 252020 17508
rect 253244 17308 253308 17372
rect 253428 17172 253492 17236
rect 221044 15948 221108 16012
rect 250852 15948 250916 16012
rect 217180 15812 217244 15876
rect 250668 15812 250732 15876
rect 218836 14724 218900 14788
rect 246804 14724 246868 14788
rect 216996 14588 217060 14652
rect 248276 14588 248340 14652
rect 211292 14452 211356 14516
rect 248092 14452 248156 14516
rect 215708 13092 215772 13156
rect 244044 13092 244108 13156
rect 214236 12956 214300 13020
rect 245516 12956 245580 13020
rect 219572 11868 219636 11932
rect 219204 11732 219268 11796
rect 242756 11732 242820 11796
rect 211108 11596 211172 11660
rect 242572 11596 242636 11660
rect 218652 10508 218716 10572
rect 237972 10508 238036 10572
rect 216628 10372 216692 10436
rect 239812 10372 239876 10436
rect 216812 10236 216876 10300
rect 239996 10236 240060 10300
rect 235580 9148 235644 9212
rect 214052 9012 214116 9076
rect 237236 9012 237300 9076
rect 209820 8876 209884 8940
rect 252140 8876 252204 8940
rect 226380 7924 226444 7988
rect 225276 7788 225340 7852
rect 223988 7652 224052 7716
rect 223804 7516 223868 7580
rect 233924 7516 233988 7580
rect 224908 6564 224972 6628
rect 3372 6428 3436 6492
rect 225092 6428 225156 6492
rect 230980 6428 231044 6492
rect 223620 6292 223684 6356
rect 233004 6292 233068 6356
rect 220860 6156 220924 6220
rect 255084 6156 255148 6220
rect 298508 5612 298572 5676
rect 229876 5340 229940 5404
rect 230060 5204 230124 5268
rect 251036 5068 251100 5132
rect 252324 4932 252388 4996
rect 253612 4796 253676 4860
rect 228956 3708 229020 3772
rect 228588 3572 228652 3636
rect 228772 3436 228836 3500
rect 249012 3436 249076 3500
rect 230244 3300 230308 3364
rect 262628 3300 262692 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 3555 446860 3621 446861
rect 3555 446796 3556 446860
rect 3620 446796 3621 446860
rect 3555 446795 3621 446796
rect 3371 446452 3437 446453
rect 3371 446388 3372 446452
rect 3436 446388 3437 446452
rect 3371 446387 3437 446388
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 6493 3434 446387
rect 3558 45525 3618 446795
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 3555 45524 3621 45525
rect 3555 45460 3556 45524
rect 3620 45460 3621 45524
rect 3555 45459 3621 45460
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 3371 6492 3437 6493
rect 3371 6428 3372 6492
rect 3436 6428 3437 6492
rect 3371 6427 3437 6428
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 691292 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 691292 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 691292 87914 700398
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 691292 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 691292 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 691292 123914 700398
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 691292 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 691292 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 691292 159914 700398
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 80952 687454 81300 687486
rect 80952 687218 81008 687454
rect 81244 687218 81300 687454
rect 80952 687134 81300 687218
rect 80952 686898 81008 687134
rect 81244 686898 81300 687134
rect 80952 686866 81300 686898
rect 169760 687454 170108 687486
rect 169760 687218 169816 687454
rect 170052 687218 170108 687454
rect 169760 687134 170108 687218
rect 169760 686898 169816 687134
rect 170052 686898 170108 687134
rect 169760 686866 170108 686898
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 80272 655954 80620 655986
rect 80272 655718 80328 655954
rect 80564 655718 80620 655954
rect 80272 655634 80620 655718
rect 80272 655398 80328 655634
rect 80564 655398 80620 655634
rect 80272 655366 80620 655398
rect 170440 655954 170788 655986
rect 170440 655718 170496 655954
rect 170732 655718 170788 655954
rect 170440 655634 170788 655718
rect 170440 655398 170496 655634
rect 170732 655398 170788 655634
rect 170440 655366 170788 655398
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 80952 651454 81300 651486
rect 80952 651218 81008 651454
rect 81244 651218 81300 651454
rect 80952 651134 81300 651218
rect 80952 650898 81008 651134
rect 81244 650898 81300 651134
rect 80952 650866 81300 650898
rect 169760 651454 170108 651486
rect 169760 651218 169816 651454
rect 170052 651218 170108 651454
rect 169760 651134 170108 651218
rect 169760 650898 169816 651134
rect 170052 650898 170108 651134
rect 169760 650866 170108 650898
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 80272 619954 80620 619986
rect 80272 619718 80328 619954
rect 80564 619718 80620 619954
rect 80272 619634 80620 619718
rect 80272 619398 80328 619634
rect 80564 619398 80620 619634
rect 80272 619366 80620 619398
rect 170440 619954 170788 619986
rect 170440 619718 170496 619954
rect 170732 619718 170788 619954
rect 170440 619634 170788 619718
rect 170440 619398 170496 619634
rect 170732 619398 170788 619634
rect 170440 619366 170788 619398
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 80952 615454 81300 615486
rect 80952 615218 81008 615454
rect 81244 615218 81300 615454
rect 80952 615134 81300 615218
rect 80952 614898 81008 615134
rect 81244 614898 81300 615134
rect 80952 614866 81300 614898
rect 169760 615454 170108 615486
rect 169760 615218 169816 615454
rect 170052 615218 170108 615454
rect 169760 615134 170108 615218
rect 169760 614898 169816 615134
rect 170052 614898 170108 615134
rect 169760 614866 170108 614898
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 92928 599450 92988 600100
rect 94288 599450 94348 600100
rect 95376 599450 95436 600100
rect 92928 599390 93042 599450
rect 92982 597413 93042 599390
rect 94270 599390 94348 599450
rect 95374 599390 95436 599450
rect 97688 599450 97748 600100
rect 98912 599450 98972 600100
rect 100000 599450 100060 600100
rect 101088 599450 101148 600100
rect 97688 599390 97826 599450
rect 92979 597412 93045 597413
rect 92979 597348 92980 597412
rect 93044 597348 93045 597412
rect 92979 597347 93045 597348
rect 94270 597005 94330 599390
rect 94267 597004 94333 597005
rect 94267 596940 94268 597004
rect 94332 596940 94333 597004
rect 94267 596939 94333 596940
rect 95374 596325 95434 599390
rect 97766 597005 97826 599390
rect 98870 599390 98972 599450
rect 99974 599390 100060 599450
rect 101078 599390 101148 599450
rect 102312 599450 102372 600100
rect 103400 599450 103460 600100
rect 104760 599450 104820 600100
rect 102312 599390 102426 599450
rect 98870 597413 98930 599390
rect 98867 597412 98933 597413
rect 98867 597348 98868 597412
rect 98932 597348 98933 597412
rect 98867 597347 98933 597348
rect 99974 597141 100034 599390
rect 101078 597413 101138 599390
rect 102366 597549 102426 599390
rect 103286 599390 103460 599450
rect 104758 599390 104820 599450
rect 105304 599450 105364 600100
rect 105712 599450 105772 600100
rect 110472 599450 110532 600100
rect 105304 599390 105370 599450
rect 102363 597548 102429 597549
rect 102363 597484 102364 597548
rect 102428 597484 102429 597548
rect 102363 597483 102429 597484
rect 101075 597412 101141 597413
rect 101075 597348 101076 597412
rect 101140 597348 101141 597412
rect 101075 597347 101141 597348
rect 103286 597277 103346 599390
rect 103283 597276 103349 597277
rect 103283 597212 103284 597276
rect 103348 597212 103349 597276
rect 103283 597211 103349 597212
rect 104758 597141 104818 599390
rect 105310 597549 105370 599390
rect 105678 599390 105772 599450
rect 110462 599390 110532 599450
rect 115504 599450 115564 600100
rect 120536 599450 120596 600100
rect 125568 599450 125628 600100
rect 115504 599390 115674 599450
rect 120536 599390 120642 599450
rect 105307 597548 105373 597549
rect 105307 597484 105308 597548
rect 105372 597484 105373 597548
rect 105307 597483 105373 597484
rect 105678 597277 105738 599390
rect 105675 597276 105741 597277
rect 105675 597212 105676 597276
rect 105740 597212 105741 597276
rect 105675 597211 105741 597212
rect 99971 597140 100037 597141
rect 99971 597076 99972 597140
rect 100036 597076 100037 597140
rect 99971 597075 100037 597076
rect 104755 597140 104821 597141
rect 104755 597076 104756 597140
rect 104820 597076 104821 597140
rect 104755 597075 104821 597076
rect 97763 597004 97829 597005
rect 97763 596940 97764 597004
rect 97828 596940 97829 597004
rect 97763 596939 97829 596940
rect 110462 596869 110522 599390
rect 110459 596868 110525 596869
rect 110459 596804 110460 596868
rect 110524 596804 110525 596868
rect 110459 596803 110525 596804
rect 115614 596325 115674 599390
rect 120582 596325 120642 599390
rect 125550 599390 125628 599450
rect 130464 599450 130524 600100
rect 135496 599450 135556 600100
rect 130464 599390 130578 599450
rect 125550 596733 125610 599390
rect 130518 597005 130578 599390
rect 135486 599390 135556 599450
rect 140528 599450 140588 600100
rect 140528 599390 140698 599450
rect 130515 597004 130581 597005
rect 130515 596940 130516 597004
rect 130580 596940 130581 597004
rect 130515 596939 130581 596940
rect 125547 596732 125613 596733
rect 125547 596668 125548 596732
rect 125612 596668 125613 596732
rect 125547 596667 125613 596668
rect 135486 596597 135546 599390
rect 140638 596597 140698 599390
rect 135483 596596 135549 596597
rect 135483 596532 135484 596596
rect 135548 596532 135549 596596
rect 135483 596531 135549 596532
rect 140635 596596 140701 596597
rect 140635 596532 140636 596596
rect 140700 596532 140701 596596
rect 140635 596531 140701 596532
rect 95371 596324 95437 596325
rect 95371 596260 95372 596324
rect 95436 596260 95437 596324
rect 95371 596259 95437 596260
rect 115611 596324 115677 596325
rect 115611 596260 115612 596324
rect 115676 596260 115677 596324
rect 115611 596259 115677 596260
rect 120579 596324 120645 596325
rect 120579 596260 120580 596324
rect 120644 596260 120645 596324
rect 120579 596259 120645 596260
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 80272 547954 80620 547986
rect 80272 547718 80328 547954
rect 80564 547718 80620 547954
rect 80272 547634 80620 547718
rect 80272 547398 80328 547634
rect 80564 547398 80620 547634
rect 80272 547366 80620 547398
rect 170440 547954 170788 547986
rect 170440 547718 170496 547954
rect 170732 547718 170788 547954
rect 170440 547634 170788 547718
rect 170440 547398 170496 547634
rect 170732 547398 170788 547634
rect 170440 547366 170788 547398
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 80952 543454 81300 543486
rect 80952 543218 81008 543454
rect 81244 543218 81300 543454
rect 80952 543134 81300 543218
rect 80952 542898 81008 543134
rect 81244 542898 81300 543134
rect 80952 542866 81300 542898
rect 169760 543454 170108 543486
rect 169760 543218 169816 543454
rect 170052 543218 170108 543454
rect 169760 543134 170108 543218
rect 169760 542898 169816 543134
rect 170052 542898 170108 543134
rect 169760 542866 170108 542898
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 80272 511954 80620 511986
rect 80272 511718 80328 511954
rect 80564 511718 80620 511954
rect 80272 511634 80620 511718
rect 80272 511398 80328 511634
rect 80564 511398 80620 511634
rect 80272 511366 80620 511398
rect 170440 511954 170788 511986
rect 170440 511718 170496 511954
rect 170732 511718 170788 511954
rect 170440 511634 170788 511718
rect 170440 511398 170496 511634
rect 170732 511398 170788 511634
rect 170440 511366 170788 511398
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 80952 507454 81300 507486
rect 80952 507218 81008 507454
rect 81244 507218 81300 507454
rect 80952 507134 81300 507218
rect 80952 506898 81008 507134
rect 81244 506898 81300 507134
rect 80952 506866 81300 506898
rect 169760 507454 170108 507486
rect 169760 507218 169816 507454
rect 170052 507218 170108 507454
rect 169760 507134 170108 507218
rect 169760 506898 169816 507134
rect 170052 506898 170108 507134
rect 169760 506866 170108 506898
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 92928 489930 92988 490106
rect 94288 489930 94348 490106
rect 95376 489930 95436 490106
rect 92928 489870 93042 489930
rect 92982 488477 93042 489870
rect 94270 489870 94348 489930
rect 95374 489870 95436 489930
rect 97688 489930 97748 490106
rect 98912 489930 98972 490106
rect 100000 489930 100060 490106
rect 101088 489930 101148 490106
rect 97688 489870 97826 489930
rect 94270 488477 94330 489870
rect 95374 488477 95434 489870
rect 97766 488477 97826 489870
rect 98870 489870 98972 489930
rect 99974 489870 100060 489930
rect 101078 489870 101148 489930
rect 102312 489930 102372 490106
rect 103400 489930 103460 490106
rect 104760 489930 104820 490106
rect 102312 489870 102426 489930
rect 98870 488477 98930 489870
rect 99974 488477 100034 489870
rect 101078 488477 101138 489870
rect 102366 488477 102426 489870
rect 103286 489870 103460 489930
rect 104758 489870 104820 489930
rect 105304 489930 105364 490106
rect 105712 489930 105772 490106
rect 110472 489930 110532 490106
rect 105304 489870 105370 489930
rect 92979 488476 93045 488477
rect 92979 488412 92980 488476
rect 93044 488412 93045 488476
rect 92979 488411 93045 488412
rect 94267 488476 94333 488477
rect 94267 488412 94268 488476
rect 94332 488412 94333 488476
rect 94267 488411 94333 488412
rect 95371 488476 95437 488477
rect 95371 488412 95372 488476
rect 95436 488412 95437 488476
rect 95371 488411 95437 488412
rect 97763 488476 97829 488477
rect 97763 488412 97764 488476
rect 97828 488412 97829 488476
rect 97763 488411 97829 488412
rect 98867 488476 98933 488477
rect 98867 488412 98868 488476
rect 98932 488412 98933 488476
rect 98867 488411 98933 488412
rect 99971 488476 100037 488477
rect 99971 488412 99972 488476
rect 100036 488412 100037 488476
rect 99971 488411 100037 488412
rect 101075 488476 101141 488477
rect 101075 488412 101076 488476
rect 101140 488412 101141 488476
rect 101075 488411 101141 488412
rect 102363 488476 102429 488477
rect 102363 488412 102364 488476
rect 102428 488412 102429 488476
rect 102363 488411 102429 488412
rect 103286 488069 103346 489870
rect 104758 488477 104818 489870
rect 104755 488476 104821 488477
rect 104755 488412 104756 488476
rect 104820 488412 104821 488476
rect 104755 488411 104821 488412
rect 105310 488205 105370 489870
rect 105678 489870 105772 489930
rect 110462 489870 110532 489930
rect 115504 489930 115564 490106
rect 120536 489930 120596 490106
rect 125568 489930 125628 490106
rect 115504 489870 115674 489930
rect 120536 489870 120642 489930
rect 105678 488477 105738 489870
rect 105675 488476 105741 488477
rect 105675 488412 105676 488476
rect 105740 488412 105741 488476
rect 105675 488411 105741 488412
rect 110462 488205 110522 489870
rect 105307 488204 105373 488205
rect 105307 488140 105308 488204
rect 105372 488140 105373 488204
rect 105307 488139 105373 488140
rect 110459 488204 110525 488205
rect 110459 488140 110460 488204
rect 110524 488140 110525 488204
rect 110459 488139 110525 488140
rect 103283 488068 103349 488069
rect 103283 488004 103284 488068
rect 103348 488004 103349 488068
rect 103283 488003 103349 488004
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 475954 78914 488000
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 480454 83414 488000
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 484954 87914 488000
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 453454 92414 488000
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 457954 96914 488000
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 462454 101414 488000
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 466954 105914 488000
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 471454 110414 488000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 475954 114914 488000
rect 115614 487253 115674 489870
rect 115611 487252 115677 487253
rect 115611 487188 115612 487252
rect 115676 487188 115677 487252
rect 115611 487187 115677 487188
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 480454 119414 488000
rect 120582 487253 120642 489870
rect 125550 489870 125628 489930
rect 130464 489930 130524 490106
rect 135496 489930 135556 490106
rect 130464 489870 130578 489930
rect 120579 487252 120645 487253
rect 120579 487188 120580 487252
rect 120644 487188 120645 487252
rect 120579 487187 120645 487188
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 484954 123914 488000
rect 125550 487253 125610 489870
rect 125547 487252 125613 487253
rect 125547 487188 125548 487252
rect 125612 487188 125613 487252
rect 125547 487187 125613 487188
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 124954 123914 160398
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 453454 128414 488000
rect 130518 487253 130578 489870
rect 135486 489870 135556 489930
rect 140528 489930 140588 490106
rect 140528 489870 140698 489930
rect 130515 487252 130581 487253
rect 130515 487188 130516 487252
rect 130580 487188 130581 487252
rect 130515 487187 130581 487188
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 457954 132914 488000
rect 135486 487253 135546 489870
rect 135483 487252 135549 487253
rect 135483 487188 135484 487252
rect 135548 487188 135549 487252
rect 135483 487187 135549 487188
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 462454 137414 488000
rect 140638 487253 140698 489870
rect 140635 487252 140701 487253
rect 140635 487188 140636 487252
rect 140700 487188 140701 487252
rect 140635 487187 140701 487188
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 466954 141914 488000
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 471454 146414 488000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 475954 150914 488000
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 480454 155414 488000
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 484954 159914 488000
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 453454 164414 488000
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 457954 168914 488000
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 462454 173414 488000
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 691292 191414 695898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 691292 195914 700398
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 691292 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 691292 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 691292 231914 700398
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 691292 258914 691398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 691292 263414 695898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 691292 267914 700398
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 190952 687454 191300 687486
rect 190952 687218 191008 687454
rect 191244 687218 191300 687454
rect 190952 687134 191300 687218
rect 190952 686898 191008 687134
rect 191244 686898 191300 687134
rect 190952 686866 191300 686898
rect 279760 687454 280108 687486
rect 279760 687218 279816 687454
rect 280052 687218 280108 687454
rect 279760 687134 280108 687218
rect 279760 686898 279816 687134
rect 280052 686898 280108 687134
rect 279760 686866 280108 686898
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 190272 655954 190620 655986
rect 190272 655718 190328 655954
rect 190564 655718 190620 655954
rect 190272 655634 190620 655718
rect 190272 655398 190328 655634
rect 190564 655398 190620 655634
rect 190272 655366 190620 655398
rect 280440 655954 280788 655986
rect 280440 655718 280496 655954
rect 280732 655718 280788 655954
rect 280440 655634 280788 655718
rect 280440 655398 280496 655634
rect 280732 655398 280788 655634
rect 280440 655366 280788 655398
rect 190952 651454 191300 651486
rect 190952 651218 191008 651454
rect 191244 651218 191300 651454
rect 190952 651134 191300 651218
rect 190952 650898 191008 651134
rect 191244 650898 191300 651134
rect 190952 650866 191300 650898
rect 279760 651454 280108 651486
rect 279760 651218 279816 651454
rect 280052 651218 280108 651454
rect 279760 651134 280108 651218
rect 279760 650898 279816 651134
rect 280052 650898 280108 651134
rect 279760 650866 280108 650898
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 190272 619954 190620 619986
rect 190272 619718 190328 619954
rect 190564 619718 190620 619954
rect 190272 619634 190620 619718
rect 190272 619398 190328 619634
rect 190564 619398 190620 619634
rect 190272 619366 190620 619398
rect 280440 619954 280788 619986
rect 280440 619718 280496 619954
rect 280732 619718 280788 619954
rect 280440 619634 280788 619718
rect 280440 619398 280496 619634
rect 280732 619398 280788 619634
rect 280440 619366 280788 619398
rect 190952 615454 191300 615486
rect 190952 615218 191008 615454
rect 191244 615218 191300 615454
rect 190952 615134 191300 615218
rect 190952 614898 191008 615134
rect 191244 614898 191300 615134
rect 190952 614866 191300 614898
rect 279760 615454 280108 615486
rect 279760 615218 279816 615454
rect 280052 615218 280108 615454
rect 279760 615134 280108 615218
rect 279760 614898 279816 615134
rect 280052 614898 280108 615134
rect 279760 614866 280108 614898
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 202928 599450 202988 600100
rect 202830 599390 202988 599450
rect 204288 599450 204348 600100
rect 205376 599450 205436 600100
rect 207688 599450 207748 600100
rect 208912 599450 208972 600100
rect 204288 599390 204362 599450
rect 205376 599390 205466 599450
rect 202830 596461 202890 599390
rect 202827 596460 202893 596461
rect 202827 596396 202828 596460
rect 202892 596396 202893 596460
rect 202827 596395 202893 596396
rect 204302 596325 204362 599390
rect 205406 597141 205466 599390
rect 207614 599390 207748 599450
rect 208902 599390 208972 599450
rect 210000 599450 210060 600100
rect 211088 599450 211148 600100
rect 212312 599450 212372 600100
rect 213400 599450 213460 600100
rect 214760 599450 214820 600100
rect 215304 599450 215364 600100
rect 215712 599450 215772 600100
rect 220472 599450 220532 600100
rect 225504 599450 225564 600100
rect 210000 599390 210066 599450
rect 211088 599390 211170 599450
rect 212312 599390 212458 599450
rect 213400 599390 213562 599450
rect 214760 599390 214850 599450
rect 215304 599390 215402 599450
rect 207614 597549 207674 599390
rect 208902 597549 208962 599390
rect 210006 597549 210066 599390
rect 211110 597549 211170 599390
rect 212398 597549 212458 599390
rect 213502 597549 213562 599390
rect 214790 597549 214850 599390
rect 215342 597549 215402 599390
rect 215710 599390 215772 599450
rect 219206 599390 220532 599450
rect 225462 599390 225564 599450
rect 230536 599450 230596 600100
rect 235568 599450 235628 600100
rect 240464 599450 240524 600100
rect 245496 599450 245556 600100
rect 250528 599450 250588 600100
rect 230536 599390 230674 599450
rect 235568 599390 235642 599450
rect 240464 599390 240610 599450
rect 245496 599390 245578 599450
rect 215710 597549 215770 599390
rect 207611 597548 207677 597549
rect 207611 597484 207612 597548
rect 207676 597484 207677 597548
rect 207611 597483 207677 597484
rect 208899 597548 208965 597549
rect 208899 597484 208900 597548
rect 208964 597484 208965 597548
rect 208899 597483 208965 597484
rect 210003 597548 210069 597549
rect 210003 597484 210004 597548
rect 210068 597484 210069 597548
rect 210003 597483 210069 597484
rect 211107 597548 211173 597549
rect 211107 597484 211108 597548
rect 211172 597484 211173 597548
rect 211107 597483 211173 597484
rect 212395 597548 212461 597549
rect 212395 597484 212396 597548
rect 212460 597484 212461 597548
rect 212395 597483 212461 597484
rect 213499 597548 213565 597549
rect 213499 597484 213500 597548
rect 213564 597484 213565 597548
rect 213499 597483 213565 597484
rect 214787 597548 214853 597549
rect 214787 597484 214788 597548
rect 214852 597484 214853 597548
rect 214787 597483 214853 597484
rect 215339 597548 215405 597549
rect 215339 597484 215340 597548
rect 215404 597484 215405 597548
rect 215339 597483 215405 597484
rect 215707 597548 215773 597549
rect 215707 597484 215708 597548
rect 215772 597484 215773 597548
rect 215707 597483 215773 597484
rect 205403 597140 205469 597141
rect 205403 597076 205404 597140
rect 205468 597076 205469 597140
rect 205403 597075 205469 597076
rect 219206 596325 219266 599390
rect 225462 597549 225522 599390
rect 225459 597548 225525 597549
rect 225459 597484 225460 597548
rect 225524 597484 225525 597548
rect 225459 597483 225525 597484
rect 230614 597277 230674 599390
rect 235582 597549 235642 599390
rect 235579 597548 235645 597549
rect 235579 597484 235580 597548
rect 235644 597484 235645 597548
rect 235579 597483 235645 597484
rect 230611 597276 230677 597277
rect 230611 597212 230612 597276
rect 230676 597212 230677 597276
rect 230611 597211 230677 597212
rect 240550 596869 240610 599390
rect 245518 597549 245578 599390
rect 250486 599390 250588 599450
rect 250486 597549 250546 599390
rect 245515 597548 245581 597549
rect 245515 597484 245516 597548
rect 245580 597484 245581 597548
rect 245515 597483 245581 597484
rect 250483 597548 250549 597549
rect 250483 597484 250484 597548
rect 250548 597484 250549 597548
rect 250483 597483 250549 597484
rect 240547 596868 240613 596869
rect 240547 596804 240548 596868
rect 240612 596804 240613 596868
rect 240547 596803 240613 596804
rect 204299 596324 204365 596325
rect 204299 596260 204300 596324
rect 204364 596260 204365 596324
rect 204299 596259 204365 596260
rect 219203 596324 219269 596325
rect 219203 596260 219204 596324
rect 219268 596260 219269 596324
rect 219203 596259 219269 596260
rect 282131 589932 282197 589933
rect 282131 589868 282132 589932
rect 282196 589868 282197 589932
rect 282131 589867 282197 589868
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 190272 547954 190620 547986
rect 190272 547718 190328 547954
rect 190564 547718 190620 547954
rect 190272 547634 190620 547718
rect 190272 547398 190328 547634
rect 190564 547398 190620 547634
rect 190272 547366 190620 547398
rect 280440 547954 280788 547986
rect 280440 547718 280496 547954
rect 280732 547718 280788 547954
rect 280440 547634 280788 547718
rect 280440 547398 280496 547634
rect 280732 547398 280788 547634
rect 280440 547366 280788 547398
rect 190952 543454 191300 543486
rect 190952 543218 191008 543454
rect 191244 543218 191300 543454
rect 190952 543134 191300 543218
rect 190952 542898 191008 543134
rect 191244 542898 191300 543134
rect 190952 542866 191300 542898
rect 279760 543454 280108 543486
rect 279760 543218 279816 543454
rect 280052 543218 280108 543454
rect 279760 543134 280108 543218
rect 279760 542898 279816 543134
rect 280052 542898 280108 543134
rect 279760 542866 280108 542898
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 190272 511954 190620 511986
rect 190272 511718 190328 511954
rect 190564 511718 190620 511954
rect 190272 511634 190620 511718
rect 190272 511398 190328 511634
rect 190564 511398 190620 511634
rect 190272 511366 190620 511398
rect 280440 511954 280788 511986
rect 280440 511718 280496 511954
rect 280732 511718 280788 511954
rect 280440 511634 280788 511718
rect 280440 511398 280496 511634
rect 280732 511398 280788 511634
rect 280440 511366 280788 511398
rect 190952 507454 191300 507486
rect 190952 507218 191008 507454
rect 191244 507218 191300 507454
rect 190952 507134 191300 507218
rect 190952 506898 191008 507134
rect 191244 506898 191300 507134
rect 190952 506866 191300 506898
rect 279760 507454 280108 507486
rect 279760 507218 279816 507454
rect 280052 507218 280108 507454
rect 279760 507134 280108 507218
rect 279760 506898 279816 507134
rect 280052 506898 280108 507134
rect 279760 506866 280108 506898
rect 202928 489930 202988 490106
rect 204288 489930 204348 490106
rect 205376 489930 205436 490106
rect 207688 489930 207748 490106
rect 208912 489930 208972 490106
rect 202928 489870 203074 489930
rect 204288 489870 204362 489930
rect 205376 489870 205466 489930
rect 203014 488205 203074 489870
rect 204302 488477 204362 489870
rect 204299 488476 204365 488477
rect 204299 488412 204300 488476
rect 204364 488412 204365 488476
rect 204299 488411 204365 488412
rect 203011 488204 203077 488205
rect 203011 488140 203012 488204
rect 203076 488140 203077 488204
rect 203011 488139 203077 488140
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 480454 191414 488000
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 484954 195914 488000
rect 203014 487253 203074 488139
rect 205406 487253 205466 489870
rect 207614 489870 207748 489930
rect 208902 489870 208972 489930
rect 210000 489930 210060 490106
rect 211088 489930 211148 490106
rect 212312 489930 212372 490106
rect 210000 489870 210066 489930
rect 211088 489870 211170 489930
rect 207614 487253 207674 489870
rect 208902 487253 208962 489870
rect 210006 487389 210066 489870
rect 211110 488341 211170 489870
rect 212214 489870 212372 489930
rect 213400 489930 213460 490106
rect 214760 489930 214820 490106
rect 215304 489930 215364 490106
rect 215712 489930 215772 490106
rect 213400 489870 213562 489930
rect 214760 489870 214850 489930
rect 215304 489870 215402 489930
rect 211107 488340 211173 488341
rect 211107 488276 211108 488340
rect 211172 488276 211173 488340
rect 211107 488275 211173 488276
rect 212214 487525 212274 489870
rect 213502 488341 213562 489870
rect 214790 488477 214850 489870
rect 214787 488476 214853 488477
rect 214787 488412 214788 488476
rect 214852 488412 214853 488476
rect 214787 488411 214853 488412
rect 213499 488340 213565 488341
rect 213499 488276 213500 488340
rect 213564 488276 213565 488340
rect 213499 488275 213565 488276
rect 212211 487524 212277 487525
rect 212211 487460 212212 487524
rect 212276 487460 212277 487524
rect 212211 487459 212277 487460
rect 210003 487388 210069 487389
rect 210003 487324 210004 487388
rect 210068 487324 210069 487388
rect 210003 487323 210069 487324
rect 215342 487253 215402 489870
rect 215710 489870 215772 489930
rect 220472 489930 220532 490106
rect 225504 489930 225564 490106
rect 220472 489870 220554 489930
rect 215710 488341 215770 489870
rect 215707 488340 215773 488341
rect 215707 488276 215708 488340
rect 215772 488276 215773 488340
rect 215707 488275 215773 488276
rect 220494 487253 220554 489870
rect 225462 489870 225564 489930
rect 230536 489930 230596 490106
rect 235568 489930 235628 490106
rect 240464 489930 240524 490106
rect 245496 489930 245556 490106
rect 250528 489930 250588 490106
rect 230536 489870 230674 489930
rect 235568 489870 235642 489930
rect 240464 489870 240610 489930
rect 245496 489870 245578 489930
rect 225462 487253 225522 489870
rect 230614 487253 230674 489870
rect 203011 487252 203077 487253
rect 203011 487188 203012 487252
rect 203076 487188 203077 487252
rect 203011 487187 203077 487188
rect 205403 487252 205469 487253
rect 205403 487188 205404 487252
rect 205468 487188 205469 487252
rect 205403 487187 205469 487188
rect 207611 487252 207677 487253
rect 207611 487188 207612 487252
rect 207676 487188 207677 487252
rect 207611 487187 207677 487188
rect 208899 487252 208965 487253
rect 208899 487188 208900 487252
rect 208964 487188 208965 487252
rect 208899 487187 208965 487188
rect 215339 487252 215405 487253
rect 215339 487188 215340 487252
rect 215404 487188 215405 487252
rect 215339 487187 215405 487188
rect 220491 487252 220557 487253
rect 220491 487188 220492 487252
rect 220556 487188 220557 487252
rect 220491 487187 220557 487188
rect 225459 487252 225525 487253
rect 225459 487188 225460 487252
rect 225524 487188 225525 487252
rect 225459 487187 225525 487188
rect 230611 487252 230677 487253
rect 230611 487188 230612 487252
rect 230676 487188 230677 487252
rect 230611 487187 230677 487188
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 231294 484954 231914 488000
rect 235582 487253 235642 489870
rect 240550 487253 240610 489870
rect 245518 487253 245578 489870
rect 250486 489870 250588 489930
rect 250486 487253 250546 489870
rect 235579 487252 235645 487253
rect 235579 487188 235580 487252
rect 235644 487188 235645 487252
rect 235579 487187 235645 487188
rect 240547 487252 240613 487253
rect 240547 487188 240548 487252
rect 240612 487188 240613 487252
rect 240547 487187 240613 487188
rect 245515 487252 245581 487253
rect 245515 487188 245516 487252
rect 245580 487188 245581 487252
rect 245515 487187 245581 487188
rect 250483 487252 250549 487253
rect 250483 487188 250484 487252
rect 250548 487188 250549 487252
rect 250483 487187 250549 487188
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 202091 446588 202157 446589
rect 202091 446524 202092 446588
rect 202156 446524 202157 446588
rect 202091 446523 202157 446524
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 381454 200414 398000
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 202094 254013 202154 446523
rect 231294 446000 231914 448398
rect 267294 484954 267914 488000
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 446000 267914 448398
rect 271794 453454 272414 488000
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 264283 445908 264349 445909
rect 264283 445844 264284 445908
rect 264348 445844 264349 445908
rect 264283 445843 264349 445844
rect 262627 445772 262693 445773
rect 262627 445708 262628 445772
rect 262692 445708 262693 445772
rect 262627 445707 262693 445708
rect 211843 444140 211909 444141
rect 211843 444076 211844 444140
rect 211908 444076 211909 444140
rect 211843 444075 211909 444076
rect 212395 444140 212461 444141
rect 212395 444076 212396 444140
rect 212460 444076 212461 444140
rect 212395 444075 212461 444076
rect 212947 444140 213013 444141
rect 212947 444076 212948 444140
rect 213012 444076 213013 444140
rect 212947 444075 213013 444076
rect 251035 444140 251101 444141
rect 251035 444076 251036 444140
rect 251100 444076 251101 444140
rect 251035 444075 251101 444076
rect 256555 444140 256621 444141
rect 256555 444076 256556 444140
rect 256620 444076 256621 444140
rect 256555 444075 256621 444076
rect 211846 442373 211906 444075
rect 211843 442372 211909 442373
rect 211843 442308 211844 442372
rect 211908 442308 211909 442372
rect 211843 442307 211909 442308
rect 212398 442237 212458 444075
rect 212950 442509 213010 444075
rect 251038 442781 251098 444075
rect 251035 442780 251101 442781
rect 251035 442716 251036 442780
rect 251100 442716 251101 442780
rect 251035 442715 251101 442716
rect 256558 442645 256618 444075
rect 256555 442644 256621 442645
rect 256555 442580 256556 442644
rect 256620 442580 256621 442644
rect 256555 442579 256621 442580
rect 212947 442508 213013 442509
rect 212947 442444 212948 442508
rect 213012 442444 213013 442508
rect 212947 442443 213013 442444
rect 212395 442236 212461 442237
rect 212395 442172 212396 442236
rect 212460 442172 212461 442236
rect 212395 442171 212461 442172
rect 219568 439954 219888 439986
rect 219568 439718 219610 439954
rect 219846 439718 219888 439954
rect 219568 439634 219888 439718
rect 219568 439398 219610 439634
rect 219846 439398 219888 439634
rect 219568 439366 219888 439398
rect 250288 439954 250608 439986
rect 250288 439718 250330 439954
rect 250566 439718 250608 439954
rect 250288 439634 250608 439718
rect 250288 439398 250330 439634
rect 250566 439398 250608 439634
rect 250288 439366 250608 439398
rect 204208 435454 204528 435486
rect 204208 435218 204250 435454
rect 204486 435218 204528 435454
rect 204208 435134 204528 435218
rect 204208 434898 204250 435134
rect 204486 434898 204528 435134
rect 204208 434866 204528 434898
rect 234928 435454 235248 435486
rect 234928 435218 234970 435454
rect 235206 435218 235248 435454
rect 234928 435134 235248 435218
rect 234928 434898 234970 435134
rect 235206 434898 235248 435134
rect 234928 434866 235248 434898
rect 219568 403954 219888 403986
rect 219568 403718 219610 403954
rect 219846 403718 219888 403954
rect 219568 403634 219888 403718
rect 219568 403398 219610 403634
rect 219846 403398 219888 403634
rect 219568 403366 219888 403398
rect 250288 403954 250608 403986
rect 250288 403718 250330 403954
rect 250566 403718 250608 403954
rect 250288 403634 250608 403718
rect 250288 403398 250330 403634
rect 250566 403398 250608 403634
rect 250288 403366 250608 403398
rect 253059 399260 253125 399261
rect 253059 399196 253060 399260
rect 253124 399196 253125 399260
rect 253059 399195 253125 399196
rect 228771 398172 228837 398173
rect 228771 398108 228772 398172
rect 228836 398108 228837 398172
rect 228771 398107 228837 398108
rect 204294 385954 204914 398000
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 202091 254012 202157 254013
rect 202091 253948 202092 254012
rect 202156 253948 202157 254012
rect 202091 253947 202157 253948
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 390454 209414 398000
rect 211107 397764 211173 397765
rect 211107 397700 211108 397764
rect 211172 397700 211173 397764
rect 211107 397699 211173 397700
rect 212763 397764 212829 397765
rect 212763 397700 212764 397764
rect 212828 397700 212829 397764
rect 212763 397699 212829 397700
rect 209819 397492 209885 397493
rect 209819 397428 209820 397492
rect 209884 397428 209885 397492
rect 209819 397427 209885 397428
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 209822 8941 209882 397427
rect 211110 11661 211170 397699
rect 211475 397628 211541 397629
rect 211475 397564 211476 397628
rect 211540 397564 211541 397628
rect 211475 397563 211541 397564
rect 211291 397492 211357 397493
rect 211291 397428 211292 397492
rect 211356 397428 211357 397492
rect 211291 397427 211357 397428
rect 211294 14517 211354 397427
rect 211478 177309 211538 397563
rect 212579 397492 212645 397493
rect 212579 397428 212580 397492
rect 212644 397428 212645 397492
rect 212579 397427 212645 397428
rect 212582 392597 212642 397427
rect 212766 395317 212826 397699
rect 212763 395316 212829 395317
rect 212763 395252 212764 395316
rect 212828 395252 212829 395316
rect 212763 395251 212829 395252
rect 213294 394954 213914 398000
rect 216627 397900 216693 397901
rect 216627 397836 216628 397900
rect 216692 397836 216693 397900
rect 216627 397835 216693 397836
rect 214419 397764 214485 397765
rect 214419 397700 214420 397764
rect 214484 397700 214485 397764
rect 214419 397699 214485 397700
rect 215339 397764 215405 397765
rect 215339 397700 215340 397764
rect 215404 397700 215405 397764
rect 215339 397699 215405 397700
rect 214051 397628 214117 397629
rect 214051 397564 214052 397628
rect 214116 397564 214117 397628
rect 214051 397563 214117 397564
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 212579 392596 212645 392597
rect 212579 392532 212580 392596
rect 212644 392532 212645 392596
rect 212579 392531 212645 392532
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 211475 177308 211541 177309
rect 211475 177244 211476 177308
rect 211540 177244 211541 177308
rect 211475 177243 211541 177244
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 211291 14516 211357 14517
rect 211291 14452 211292 14516
rect 211356 14452 211357 14516
rect 211291 14451 211357 14452
rect 211107 11660 211173 11661
rect 211107 11596 211108 11660
rect 211172 11596 211173 11660
rect 211107 11595 211173 11596
rect 209819 8940 209885 8941
rect 209819 8876 209820 8940
rect 209884 8876 209885 8940
rect 209819 8875 209885 8876
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 -7066 213914 34398
rect 214054 9077 214114 397563
rect 214235 397492 214301 397493
rect 214235 397428 214236 397492
rect 214300 397428 214301 397492
rect 214235 397427 214301 397428
rect 214238 13021 214298 397427
rect 214422 177445 214482 397699
rect 215342 395589 215402 397699
rect 215707 397628 215773 397629
rect 215707 397564 215708 397628
rect 215772 397564 215773 397628
rect 215707 397563 215773 397564
rect 215523 397492 215589 397493
rect 215523 397428 215524 397492
rect 215588 397428 215589 397492
rect 215523 397427 215589 397428
rect 215339 395588 215405 395589
rect 215339 395524 215340 395588
rect 215404 395524 215405 395588
rect 215339 395523 215405 395524
rect 215526 177581 215586 397427
rect 215523 177580 215589 177581
rect 215523 177516 215524 177580
rect 215588 177516 215589 177580
rect 215523 177515 215589 177516
rect 214419 177444 214485 177445
rect 214419 177380 214420 177444
rect 214484 177380 214485 177444
rect 214419 177379 214485 177380
rect 215710 13157 215770 397563
rect 215707 13156 215773 13157
rect 215707 13092 215708 13156
rect 215772 13092 215773 13156
rect 215707 13091 215773 13092
rect 214235 13020 214301 13021
rect 214235 12956 214236 13020
rect 214300 12956 214301 13020
rect 214235 12955 214301 12956
rect 216630 10437 216690 397835
rect 217179 397764 217245 397765
rect 217179 397700 217180 397764
rect 217244 397700 217245 397764
rect 217179 397699 217245 397700
rect 216995 397628 217061 397629
rect 216995 397564 216996 397628
rect 217060 397564 217061 397628
rect 216995 397563 217061 397564
rect 216811 397492 216877 397493
rect 216811 397428 216812 397492
rect 216876 397428 216877 397492
rect 216811 397427 216877 397428
rect 216627 10436 216693 10437
rect 216627 10372 216628 10436
rect 216692 10372 216693 10436
rect 216627 10371 216693 10372
rect 216814 10301 216874 397427
rect 216998 14653 217058 397563
rect 217182 15877 217242 397699
rect 217794 363454 218414 398000
rect 219019 397764 219085 397765
rect 219019 397700 219020 397764
rect 219084 397700 219085 397764
rect 219019 397699 219085 397700
rect 221227 397764 221293 397765
rect 221227 397700 221228 397764
rect 221292 397700 221293 397764
rect 221227 397699 221293 397700
rect 222147 397764 222213 397765
rect 222147 397700 222148 397764
rect 222212 397700 222213 397764
rect 222147 397699 222213 397700
rect 218835 397628 218901 397629
rect 218835 397564 218836 397628
rect 218900 397564 218901 397628
rect 218835 397563 218901 397564
rect 218651 397492 218717 397493
rect 218651 397428 218652 397492
rect 218716 397428 218717 397492
rect 218651 397427 218717 397428
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217179 15876 217245 15877
rect 217179 15812 217180 15876
rect 217244 15812 217245 15876
rect 217179 15811 217245 15812
rect 216995 14652 217061 14653
rect 216995 14588 216996 14652
rect 217060 14588 217061 14652
rect 216995 14587 217061 14588
rect 216811 10300 216877 10301
rect 216811 10236 216812 10300
rect 216876 10236 216877 10300
rect 216811 10235 216877 10236
rect 214051 9076 214117 9077
rect 214051 9012 214052 9076
rect 214116 9012 214117 9076
rect 214051 9011 214117 9012
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 3454 218414 38898
rect 218654 10573 218714 397427
rect 218838 14789 218898 397563
rect 219022 355333 219082 397699
rect 219571 397628 219637 397629
rect 219571 397564 219572 397628
rect 219636 397564 219637 397628
rect 219571 397563 219637 397564
rect 220859 397628 220925 397629
rect 220859 397564 220860 397628
rect 220924 397564 220925 397628
rect 220859 397563 220925 397564
rect 219387 397492 219453 397493
rect 219387 397428 219388 397492
rect 219452 397428 219453 397492
rect 219387 397427 219453 397428
rect 219390 389190 219450 397427
rect 219206 389130 219450 389190
rect 219019 355332 219085 355333
rect 219019 355268 219020 355332
rect 219084 355268 219085 355332
rect 219019 355267 219085 355268
rect 218835 14788 218901 14789
rect 218835 14724 218836 14788
rect 218900 14724 218901 14788
rect 218835 14723 218901 14724
rect 219206 11797 219266 389130
rect 219574 11933 219634 397563
rect 219755 397492 219821 397493
rect 219755 397428 219756 397492
rect 219820 397428 219821 397492
rect 219755 397427 219821 397428
rect 219758 177717 219818 397427
rect 219755 177716 219821 177717
rect 219755 177652 219756 177716
rect 219820 177652 219821 177716
rect 219755 177651 219821 177652
rect 219571 11932 219637 11933
rect 219571 11868 219572 11932
rect 219636 11868 219637 11932
rect 219571 11867 219637 11868
rect 219203 11796 219269 11797
rect 219203 11732 219204 11796
rect 219268 11732 219269 11796
rect 219203 11731 219269 11732
rect 218651 10572 218717 10573
rect 218651 10508 218652 10572
rect 218716 10508 218717 10572
rect 218651 10507 218717 10508
rect 220862 6221 220922 397563
rect 221043 397492 221109 397493
rect 221043 397428 221044 397492
rect 221108 397428 221109 397492
rect 221043 397427 221109 397428
rect 221046 16013 221106 397427
rect 221230 394773 221290 397699
rect 221411 397628 221477 397629
rect 221411 397564 221412 397628
rect 221476 397564 221477 397628
rect 221411 397563 221477 397564
rect 221227 394772 221293 394773
rect 221227 394708 221228 394772
rect 221292 394708 221293 394772
rect 221227 394707 221293 394708
rect 221414 393957 221474 397563
rect 222150 396949 222210 397699
rect 222147 396948 222213 396949
rect 222147 396884 222148 396948
rect 222212 396884 222213 396948
rect 222147 396883 222213 396884
rect 221411 393956 221477 393957
rect 221411 393892 221412 393956
rect 221476 393892 221477 393956
rect 221411 393891 221477 393892
rect 222294 367954 222914 398000
rect 225459 397900 225525 397901
rect 225459 397836 225460 397900
rect 225524 397836 225525 397900
rect 225459 397835 225525 397836
rect 223803 397764 223869 397765
rect 223803 397700 223804 397764
rect 223868 397700 223869 397764
rect 223803 397699 223869 397700
rect 224907 397764 224973 397765
rect 224907 397700 224908 397764
rect 224972 397700 224973 397764
rect 224907 397699 224973 397700
rect 223067 397492 223133 397493
rect 223067 397428 223068 397492
rect 223132 397428 223133 397492
rect 223067 397427 223133 397428
rect 223619 397492 223685 397493
rect 223619 397428 223620 397492
rect 223684 397428 223685 397492
rect 223619 397427 223685 397428
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 223070 352613 223130 397427
rect 223067 352612 223133 352613
rect 223067 352548 223068 352612
rect 223132 352548 223133 352612
rect 223067 352547 223133 352548
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 221043 16012 221109 16013
rect 221043 15948 221044 16012
rect 221108 15948 221109 16012
rect 221043 15947 221109 15948
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 220859 6220 220925 6221
rect 220859 6156 220860 6220
rect 220924 6156 220925 6220
rect 220859 6155 220925 6156
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 -1306 222914 7398
rect 223622 6357 223682 397427
rect 223806 7581 223866 397699
rect 223987 397628 224053 397629
rect 223987 397564 223988 397628
rect 224052 397564 224053 397628
rect 224910 397626 224970 397699
rect 223987 397563 224053 397564
rect 224726 397566 224970 397626
rect 225091 397628 225157 397629
rect 223990 7717 224050 397563
rect 224171 397492 224237 397493
rect 224171 397428 224172 397492
rect 224236 397428 224237 397492
rect 224171 397427 224237 397428
rect 224174 351117 224234 397427
rect 224726 389190 224786 397566
rect 225091 397564 225092 397628
rect 225156 397564 225157 397628
rect 225091 397563 225157 397564
rect 224726 389130 224970 389190
rect 224171 351116 224237 351117
rect 224171 351052 224172 351116
rect 224236 351052 224237 351116
rect 224171 351051 224237 351052
rect 223987 7716 224053 7717
rect 223987 7652 223988 7716
rect 224052 7652 224053 7716
rect 223987 7651 224053 7652
rect 223803 7580 223869 7581
rect 223803 7516 223804 7580
rect 223868 7516 223869 7580
rect 223803 7515 223869 7516
rect 224910 6629 224970 389130
rect 224907 6628 224973 6629
rect 224907 6564 224908 6628
rect 224972 6564 224973 6628
rect 224907 6563 224973 6564
rect 225094 6493 225154 397563
rect 225275 397492 225341 397493
rect 225275 397428 225276 397492
rect 225340 397428 225341 397492
rect 225275 397427 225341 397428
rect 225278 7853 225338 397427
rect 225462 392733 225522 397835
rect 226563 397628 226629 397629
rect 226563 397564 226564 397628
rect 226628 397564 226629 397628
rect 226563 397563 226629 397564
rect 226379 397492 226445 397493
rect 226379 397428 226380 397492
rect 226444 397428 226445 397492
rect 226379 397427 226445 397428
rect 225459 392732 225525 392733
rect 225459 392668 225460 392732
rect 225524 392668 225525 392732
rect 225459 392667 225525 392668
rect 226382 7989 226442 397427
rect 226566 392869 226626 397563
rect 226563 392868 226629 392869
rect 226563 392804 226564 392868
rect 226628 392804 226629 392868
rect 226563 392803 226629 392804
rect 226794 372454 227414 398000
rect 228587 397628 228653 397629
rect 228587 397564 228588 397628
rect 228652 397564 228653 397628
rect 228587 397563 228653 397564
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226379 7988 226445 7989
rect 226379 7924 226380 7988
rect 226444 7924 226445 7988
rect 226379 7923 226445 7924
rect 225275 7852 225341 7853
rect 225275 7788 225276 7852
rect 225340 7788 225341 7852
rect 225275 7787 225341 7788
rect 225091 6492 225157 6493
rect 225091 6428 225092 6492
rect 225156 6428 225157 6492
rect 225091 6427 225157 6428
rect 223619 6356 223685 6357
rect 223619 6292 223620 6356
rect 223684 6292 223685 6356
rect 223619 6291 223685 6292
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 -2266 227414 11898
rect 228590 3637 228650 397563
rect 228587 3636 228653 3637
rect 228587 3572 228588 3636
rect 228652 3572 228653 3636
rect 228587 3571 228653 3572
rect 228774 3501 228834 398107
rect 230427 397900 230493 397901
rect 230427 397836 230428 397900
rect 230492 397836 230493 397900
rect 230427 397835 230493 397836
rect 229875 397764 229941 397765
rect 229875 397700 229876 397764
rect 229940 397700 229941 397764
rect 229875 397699 229941 397700
rect 228955 397492 229021 397493
rect 228955 397428 228956 397492
rect 229020 397428 229021 397492
rect 228955 397427 229021 397428
rect 228958 3773 229018 397427
rect 229878 5405 229938 397699
rect 230059 397628 230125 397629
rect 230059 397564 230060 397628
rect 230124 397564 230125 397628
rect 230059 397563 230125 397564
rect 229875 5404 229941 5405
rect 229875 5340 229876 5404
rect 229940 5340 229941 5404
rect 229875 5339 229941 5340
rect 230062 5269 230122 397563
rect 230243 397492 230309 397493
rect 230243 397428 230244 397492
rect 230308 397428 230309 397492
rect 230243 397427 230309 397428
rect 230059 5268 230125 5269
rect 230059 5204 230060 5268
rect 230124 5204 230125 5268
rect 230059 5203 230125 5204
rect 228955 3772 229021 3773
rect 228955 3708 228956 3772
rect 229020 3708 229021 3772
rect 228955 3707 229021 3708
rect 228771 3500 228837 3501
rect 228771 3436 228772 3500
rect 228836 3436 228837 3500
rect 228771 3435 228837 3436
rect 230246 3365 230306 397427
rect 230430 395453 230490 397835
rect 230611 397764 230677 397765
rect 230611 397700 230612 397764
rect 230676 397700 230677 397764
rect 230611 397699 230677 397700
rect 230427 395452 230493 395453
rect 230427 395388 230428 395452
rect 230492 395388 230493 395452
rect 230427 395387 230493 395388
rect 230614 177309 230674 397699
rect 230795 397628 230861 397629
rect 230795 397564 230796 397628
rect 230860 397564 230861 397628
rect 230795 397563 230861 397564
rect 230611 177308 230677 177309
rect 230611 177244 230612 177308
rect 230676 177244 230677 177308
rect 230611 177243 230677 177244
rect 230798 18597 230858 397563
rect 230979 397492 231045 397493
rect 230979 397428 230980 397492
rect 231044 397428 231045 397492
rect 230979 397427 231045 397428
rect 230795 18596 230861 18597
rect 230795 18532 230796 18596
rect 230860 18532 230861 18596
rect 230795 18531 230861 18532
rect 230982 6493 231042 397427
rect 231294 376954 231914 398000
rect 233187 397900 233253 397901
rect 233187 397836 233188 397900
rect 233252 397836 233253 397900
rect 233187 397835 233253 397836
rect 232635 397764 232701 397765
rect 232635 397700 232636 397764
rect 232700 397700 232701 397764
rect 232635 397699 232701 397700
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 232638 20093 232698 397699
rect 232819 397628 232885 397629
rect 232819 397564 232820 397628
rect 232884 397564 232885 397628
rect 232819 397563 232885 397564
rect 232822 20229 232882 397563
rect 233003 397492 233069 397493
rect 233003 397428 233004 397492
rect 233068 397428 233069 397492
rect 233003 397427 233069 397428
rect 232819 20228 232885 20229
rect 232819 20164 232820 20228
rect 232884 20164 232885 20228
rect 232819 20163 232885 20164
rect 232635 20092 232701 20093
rect 232635 20028 232636 20092
rect 232700 20028 232701 20092
rect 232635 20027 232701 20028
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 230979 6492 231045 6493
rect 230979 6428 230980 6492
rect 231044 6428 231045 6492
rect 230979 6427 231045 6428
rect 230243 3364 230309 3365
rect 230243 3300 230244 3364
rect 230308 3300 230309 3364
rect 230243 3299 230309 3300
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 -3226 231914 16398
rect 233006 6357 233066 397427
rect 233190 393957 233250 397835
rect 233923 397764 233989 397765
rect 233923 397700 233924 397764
rect 233988 397700 233989 397764
rect 233923 397699 233989 397700
rect 235211 397764 235277 397765
rect 235211 397700 235212 397764
rect 235276 397700 235277 397764
rect 235211 397699 235277 397700
rect 233187 393956 233253 393957
rect 233187 393892 233188 393956
rect 233252 393892 233253 393956
rect 233187 393891 233253 393892
rect 233926 7581 233986 397699
rect 234107 397628 234173 397629
rect 234107 397564 234108 397628
rect 234172 397564 234173 397628
rect 234107 397563 234173 397564
rect 234110 86325 234170 397563
rect 234291 397492 234357 397493
rect 234291 397428 234292 397492
rect 234356 397428 234357 397492
rect 234291 397427 234357 397428
rect 234107 86324 234173 86325
rect 234107 86260 234108 86324
rect 234172 86260 234173 86324
rect 234107 86259 234173 86260
rect 234294 19957 234354 397427
rect 235214 355333 235274 397699
rect 235395 397628 235461 397629
rect 235395 397564 235396 397628
rect 235460 397564 235461 397628
rect 235395 397563 235461 397564
rect 235211 355332 235277 355333
rect 235211 355268 235212 355332
rect 235276 355268 235277 355332
rect 235211 355267 235277 355268
rect 235398 25669 235458 397563
rect 235579 397492 235645 397493
rect 235579 397428 235580 397492
rect 235644 397428 235645 397492
rect 235579 397427 235645 397428
rect 235395 25668 235461 25669
rect 235395 25604 235396 25668
rect 235460 25604 235461 25668
rect 235395 25603 235461 25604
rect 234291 19956 234357 19957
rect 234291 19892 234292 19956
rect 234356 19892 234357 19956
rect 234291 19891 234357 19892
rect 235582 9213 235642 397427
rect 235794 381454 236414 398000
rect 236867 397764 236933 397765
rect 236867 397700 236868 397764
rect 236932 397700 236933 397764
rect 236867 397699 236933 397700
rect 237971 397764 238037 397765
rect 237971 397700 237972 397764
rect 238036 397700 238037 397764
rect 237971 397699 238037 397700
rect 239443 397764 239509 397765
rect 239443 397700 239444 397764
rect 239508 397700 239509 397764
rect 239443 397699 239509 397700
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 236870 84829 236930 397699
rect 237051 397628 237117 397629
rect 237051 397564 237052 397628
rect 237116 397564 237117 397628
rect 237051 397563 237117 397564
rect 236867 84828 236933 84829
rect 236867 84764 236868 84828
rect 236932 84764 236933 84828
rect 236867 84763 236933 84764
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 237054 21589 237114 397563
rect 237235 397492 237301 397493
rect 237235 397428 237236 397492
rect 237300 397428 237301 397492
rect 237235 397427 237301 397428
rect 237051 21588 237117 21589
rect 237051 21524 237052 21588
rect 237116 21524 237117 21588
rect 237051 21523 237117 21524
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235579 9212 235645 9213
rect 235579 9148 235580 9212
rect 235644 9148 235645 9212
rect 235579 9147 235645 9148
rect 233923 7580 233989 7581
rect 233923 7516 233924 7580
rect 233988 7516 233989 7580
rect 233923 7515 233989 7516
rect 233003 6356 233069 6357
rect 233003 6292 233004 6356
rect 233068 6292 233069 6356
rect 233003 6291 233069 6292
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 -4186 236414 20898
rect 237238 9077 237298 397427
rect 237974 10573 238034 397699
rect 238155 397628 238221 397629
rect 238155 397564 238156 397628
rect 238220 397564 238221 397628
rect 238155 397563 238221 397564
rect 238158 354109 238218 397563
rect 238339 397492 238405 397493
rect 238339 397428 238340 397492
rect 238404 397428 238405 397492
rect 238339 397427 238405 397428
rect 238155 354108 238221 354109
rect 238155 354044 238156 354108
rect 238220 354044 238221 354108
rect 238155 354043 238221 354044
rect 238342 21453 238402 397427
rect 239446 22949 239506 397699
rect 239627 397628 239693 397629
rect 239627 397564 239628 397628
rect 239692 397564 239693 397628
rect 239627 397563 239693 397564
rect 239443 22948 239509 22949
rect 239443 22884 239444 22948
rect 239508 22884 239509 22948
rect 239443 22883 239509 22884
rect 238339 21452 238405 21453
rect 238339 21388 238340 21452
rect 238404 21388 238405 21452
rect 238339 21387 238405 21388
rect 239630 21317 239690 397563
rect 239811 397492 239877 397493
rect 239811 397428 239812 397492
rect 239876 397428 239877 397492
rect 239811 397427 239877 397428
rect 239995 397492 240061 397493
rect 239995 397428 239996 397492
rect 240060 397428 240061 397492
rect 239995 397427 240061 397428
rect 239627 21316 239693 21317
rect 239627 21252 239628 21316
rect 239692 21252 239693 21316
rect 239627 21251 239693 21252
rect 237971 10572 238037 10573
rect 237971 10508 237972 10572
rect 238036 10508 238037 10572
rect 237971 10507 238037 10508
rect 239814 10437 239874 397427
rect 239811 10436 239877 10437
rect 239811 10372 239812 10436
rect 239876 10372 239877 10436
rect 239811 10371 239877 10372
rect 239998 10301 240058 397427
rect 240294 385954 240914 398000
rect 242387 397900 242453 397901
rect 242387 397836 242388 397900
rect 242452 397836 242453 397900
rect 242387 397835 242453 397836
rect 242203 397764 242269 397765
rect 242203 397700 242204 397764
rect 242268 397700 242269 397764
rect 242203 397699 242269 397700
rect 241099 397492 241165 397493
rect 241099 397428 241100 397492
rect 241164 397428 241165 397492
rect 241099 397427 241165 397428
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 241102 82109 241162 397427
rect 241099 82108 241165 82109
rect 241099 82044 241100 82108
rect 241164 82044 241165 82108
rect 241099 82043 241165 82044
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 239995 10300 240061 10301
rect 239995 10236 239996 10300
rect 240060 10236 240061 10300
rect 239995 10235 240061 10236
rect 237235 9076 237301 9077
rect 237235 9012 237236 9076
rect 237300 9012 237301 9076
rect 237235 9011 237301 9012
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 -5146 240914 25398
rect 242206 22813 242266 397699
rect 242203 22812 242269 22813
rect 242203 22748 242204 22812
rect 242268 22748 242269 22812
rect 242203 22747 242269 22748
rect 242390 22677 242450 397835
rect 243675 397764 243741 397765
rect 243675 397700 243676 397764
rect 243740 397700 243741 397764
rect 243675 397699 243741 397700
rect 242755 397628 242821 397629
rect 242755 397564 242756 397628
rect 242820 397564 242821 397628
rect 242755 397563 242821 397564
rect 242571 397492 242637 397493
rect 242571 397428 242572 397492
rect 242636 397428 242637 397492
rect 242571 397427 242637 397428
rect 242387 22676 242453 22677
rect 242387 22612 242388 22676
rect 242452 22612 242453 22676
rect 242387 22611 242453 22612
rect 242574 11661 242634 397427
rect 242758 11797 242818 397563
rect 243678 352885 243738 397699
rect 243859 397628 243925 397629
rect 243859 397564 243860 397628
rect 243924 397564 243925 397628
rect 243859 397563 243925 397564
rect 243675 352884 243741 352885
rect 243675 352820 243676 352884
rect 243740 352820 243741 352884
rect 243675 352819 243741 352820
rect 243862 24445 243922 397563
rect 244043 397492 244109 397493
rect 244043 397428 244044 397492
rect 244108 397428 244109 397492
rect 244043 397427 244109 397428
rect 243859 24444 243925 24445
rect 243859 24380 243860 24444
rect 243924 24380 243925 24444
rect 243859 24379 243925 24380
rect 244046 13157 244106 397427
rect 244794 390454 245414 398000
rect 246987 397900 247053 397901
rect 246987 397836 246988 397900
rect 247052 397836 247053 397900
rect 246987 397835 247053 397836
rect 247723 397900 247789 397901
rect 247723 397836 247724 397900
rect 247788 397836 247789 397900
rect 247723 397835 247789 397836
rect 246619 397764 246685 397765
rect 246619 397700 246620 397764
rect 246684 397700 246685 397764
rect 246619 397699 246685 397700
rect 246435 397628 246501 397629
rect 246435 397564 246436 397628
rect 246500 397564 246501 397628
rect 246435 397563 246501 397564
rect 245515 397492 245581 397493
rect 245515 397428 245516 397492
rect 245580 397428 245581 397492
rect 245515 397427 245581 397428
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244043 13156 244109 13157
rect 244043 13092 244044 13156
rect 244108 13092 244109 13156
rect 244043 13091 244109 13092
rect 242755 11796 242821 11797
rect 242755 11732 242756 11796
rect 242820 11732 242821 11796
rect 242755 11731 242821 11732
rect 242571 11660 242637 11661
rect 242571 11596 242572 11660
rect 242636 11596 242637 11660
rect 242571 11595 242637 11596
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 -6106 245414 29898
rect 245518 13021 245578 397427
rect 246438 24309 246498 397563
rect 246435 24308 246501 24309
rect 246435 24244 246436 24308
rect 246500 24244 246501 24308
rect 246435 24243 246501 24244
rect 246622 24173 246682 397699
rect 246803 397492 246869 397493
rect 246803 397428 246804 397492
rect 246868 397428 246869 397492
rect 246803 397427 246869 397428
rect 246619 24172 246685 24173
rect 246619 24108 246620 24172
rect 246684 24108 246685 24172
rect 246619 24107 246685 24108
rect 246806 14789 246866 397427
rect 246990 395589 247050 397835
rect 246987 395588 247053 395589
rect 246987 395524 246988 395588
rect 247052 395524 247053 395588
rect 246987 395523 247053 395524
rect 247726 352749 247786 397835
rect 247907 397764 247973 397765
rect 247907 397700 247908 397764
rect 247972 397700 247973 397764
rect 247907 397699 247973 397700
rect 248643 397764 248709 397765
rect 248643 397700 248644 397764
rect 248708 397700 248709 397764
rect 248643 397699 248709 397700
rect 247723 352748 247789 352749
rect 247723 352684 247724 352748
rect 247788 352684 247789 352748
rect 247723 352683 247789 352684
rect 247910 26893 247970 397699
rect 248091 397628 248157 397629
rect 248091 397564 248092 397628
rect 248156 397564 248157 397628
rect 248091 397563 248157 397564
rect 247907 26892 247973 26893
rect 247907 26828 247908 26892
rect 247972 26828 247973 26892
rect 247907 26827 247973 26828
rect 246803 14788 246869 14789
rect 246803 14724 246804 14788
rect 246868 14724 246869 14788
rect 246803 14723 246869 14724
rect 248094 14517 248154 397563
rect 248275 397492 248341 397493
rect 248275 397428 248276 397492
rect 248340 397428 248341 397492
rect 248275 397427 248341 397428
rect 248278 14653 248338 397427
rect 248646 352613 248706 397699
rect 248827 397628 248893 397629
rect 248827 397564 248828 397628
rect 248892 397564 248893 397628
rect 248827 397563 248893 397564
rect 248643 352612 248709 352613
rect 248643 352548 248644 352612
rect 248708 352548 248709 352612
rect 248643 352547 248709 352548
rect 248830 86189 248890 397563
rect 249011 397492 249077 397493
rect 249011 397428 249012 397492
rect 249076 397428 249077 397492
rect 249011 397427 249077 397428
rect 248827 86188 248893 86189
rect 248827 86124 248828 86188
rect 248892 86124 248893 86188
rect 248827 86123 248893 86124
rect 248275 14652 248341 14653
rect 248275 14588 248276 14652
rect 248340 14588 248341 14652
rect 248275 14587 248341 14588
rect 248091 14516 248157 14517
rect 248091 14452 248092 14516
rect 248156 14452 248157 14516
rect 248091 14451 248157 14452
rect 245515 13020 245581 13021
rect 245515 12956 245516 13020
rect 245580 12956 245581 13020
rect 245515 12955 245581 12956
rect 249014 3501 249074 397427
rect 249294 394954 249914 398000
rect 251955 397900 252021 397901
rect 251955 397836 251956 397900
rect 252020 397836 252021 397900
rect 251955 397835 252021 397836
rect 250667 397764 250733 397765
rect 250667 397700 250668 397764
rect 250732 397700 250733 397764
rect 250667 397699 250733 397700
rect 251771 397764 251837 397765
rect 251771 397700 251772 397764
rect 251836 397700 251837 397764
rect 251771 397699 251837 397700
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249011 3500 249077 3501
rect 249011 3436 249012 3500
rect 249076 3436 249077 3500
rect 249011 3435 249077 3436
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 -7066 249914 34398
rect 250670 15877 250730 397699
rect 250851 397628 250917 397629
rect 250851 397564 250852 397628
rect 250916 397564 250917 397628
rect 250851 397563 250917 397564
rect 250854 16013 250914 397563
rect 251035 397492 251101 397493
rect 251035 397428 251036 397492
rect 251100 397428 251101 397492
rect 251035 397427 251101 397428
rect 250851 16012 250917 16013
rect 250851 15948 250852 16012
rect 250916 15948 250917 16012
rect 250851 15947 250917 15948
rect 250667 15876 250733 15877
rect 250667 15812 250668 15876
rect 250732 15812 250733 15876
rect 250667 15811 250733 15812
rect 251038 5133 251098 397427
rect 251774 353973 251834 397699
rect 251771 353972 251837 353973
rect 251771 353908 251772 353972
rect 251836 353908 251837 353972
rect 251771 353907 251837 353908
rect 251958 17509 252018 397835
rect 252139 397628 252205 397629
rect 252139 397564 252140 397628
rect 252204 397564 252205 397628
rect 252139 397563 252205 397564
rect 251955 17508 252021 17509
rect 251955 17444 251956 17508
rect 252020 17444 252021 17508
rect 251955 17443 252021 17444
rect 252142 8941 252202 397563
rect 252323 397492 252389 397493
rect 252323 397428 252324 397492
rect 252388 397428 252389 397492
rect 252323 397427 252389 397428
rect 252139 8940 252205 8941
rect 252139 8876 252140 8940
rect 252204 8876 252205 8940
rect 252139 8875 252205 8876
rect 251035 5132 251101 5133
rect 251035 5068 251036 5132
rect 251100 5068 251101 5132
rect 251035 5067 251101 5068
rect 252326 4997 252386 397427
rect 253062 395317 253122 399195
rect 254531 398852 254597 398853
rect 254531 398788 254532 398852
rect 254596 398788 254597 398852
rect 254531 398787 254597 398788
rect 253427 397764 253493 397765
rect 253427 397700 253428 397764
rect 253492 397700 253493 397764
rect 253427 397699 253493 397700
rect 253243 397628 253309 397629
rect 253243 397564 253244 397628
rect 253308 397564 253309 397628
rect 253243 397563 253309 397564
rect 253059 395316 253125 395317
rect 253059 395252 253060 395316
rect 253124 395252 253125 395316
rect 253059 395251 253125 395252
rect 253246 17373 253306 397563
rect 253243 17372 253309 17373
rect 253243 17308 253244 17372
rect 253308 17308 253309 17372
rect 253243 17307 253309 17308
rect 253430 17237 253490 397699
rect 253611 397492 253677 397493
rect 253611 397428 253612 397492
rect 253676 397428 253677 397492
rect 253611 397427 253677 397428
rect 253427 17236 253493 17237
rect 253427 17172 253428 17236
rect 253492 17172 253493 17236
rect 253427 17171 253493 17172
rect 252323 4996 252389 4997
rect 252323 4932 252324 4996
rect 252388 4932 252389 4996
rect 252323 4931 252389 4932
rect 253614 4861 253674 397427
rect 253794 363454 254414 398000
rect 254534 397901 254594 398787
rect 254531 397900 254597 397901
rect 254531 397836 254532 397900
rect 254596 397836 254597 397900
rect 254531 397835 254597 397836
rect 254715 397764 254781 397765
rect 254715 397700 254716 397764
rect 254780 397700 254781 397764
rect 254715 397699 254781 397700
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 254718 87549 254778 397699
rect 254899 397628 254965 397629
rect 254899 397564 254900 397628
rect 254964 397564 254965 397628
rect 254899 397563 254965 397564
rect 254715 87548 254781 87549
rect 254715 87484 254716 87548
rect 254780 87484 254781 87548
rect 254715 87483 254781 87484
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253611 4860 253677 4861
rect 253611 4796 253612 4860
rect 253676 4796 253677 4860
rect 253611 4795 253677 4796
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3454 254414 38898
rect 254902 25533 254962 397563
rect 255083 397492 255149 397493
rect 255083 397428 255084 397492
rect 255148 397428 255149 397492
rect 255083 397427 255149 397428
rect 254899 25532 254965 25533
rect 254899 25468 254900 25532
rect 254964 25468 254965 25532
rect 254899 25467 254965 25468
rect 255086 6221 255146 397427
rect 258294 367954 258914 398000
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 255083 6220 255149 6221
rect 255083 6156 255084 6220
rect 255148 6156 255149 6220
rect 255083 6155 255149 6156
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 -1306 258914 7398
rect 262630 3365 262690 445707
rect 262811 445092 262877 445093
rect 262811 445028 262812 445092
rect 262876 445028 262877 445092
rect 262811 445027 262877 445028
rect 262814 398717 262874 445027
rect 264099 443596 264165 443597
rect 264099 443532 264100 443596
rect 264164 443532 264165 443596
rect 264099 443531 264165 443532
rect 262811 398716 262877 398717
rect 262811 398652 262812 398716
rect 262876 398652 262877 398716
rect 262811 398651 262877 398652
rect 262794 372454 263414 398000
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 264102 31789 264162 443531
rect 264286 398853 264346 445843
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 264283 398852 264349 398853
rect 264283 398788 264284 398852
rect 264348 398788 264349 398852
rect 264283 398787 264349 398788
rect 267294 376954 267914 398000
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 264099 31788 264165 31789
rect 264099 31724 264100 31788
rect 264164 31724 264165 31788
rect 264099 31723 264165 31724
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262627 3364 262693 3365
rect 262627 3300 262628 3364
rect 262692 3300 262693 3364
rect 262627 3299 262693 3300
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 457954 276914 488000
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 462454 281414 488000
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 282134 446453 282194 589867
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 282131 446452 282197 446453
rect 282131 446388 282132 446452
rect 282196 446388 282197 446452
rect 282131 446387 282197 446388
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 691292 299414 695898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 691292 303914 700398
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 691292 330914 691398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 691292 335414 695898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 691292 339914 700398
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 691292 366914 691398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 691292 371414 695898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 691292 375914 700398
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 300952 687454 301300 687486
rect 300952 687218 301008 687454
rect 301244 687218 301300 687454
rect 300952 687134 301300 687218
rect 300952 686898 301008 687134
rect 301244 686898 301300 687134
rect 300952 686866 301300 686898
rect 389760 687454 390108 687486
rect 389760 687218 389816 687454
rect 390052 687218 390108 687454
rect 389760 687134 390108 687218
rect 389760 686898 389816 687134
rect 390052 686898 390108 687134
rect 389760 686866 390108 686898
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 300272 655954 300620 655986
rect 300272 655718 300328 655954
rect 300564 655718 300620 655954
rect 300272 655634 300620 655718
rect 300272 655398 300328 655634
rect 300564 655398 300620 655634
rect 300272 655366 300620 655398
rect 390440 655954 390788 655986
rect 390440 655718 390496 655954
rect 390732 655718 390788 655954
rect 390440 655634 390788 655718
rect 390440 655398 390496 655634
rect 390732 655398 390788 655634
rect 390440 655366 390788 655398
rect 300952 651454 301300 651486
rect 300952 651218 301008 651454
rect 301244 651218 301300 651454
rect 300952 651134 301300 651218
rect 300952 650898 301008 651134
rect 301244 650898 301300 651134
rect 300952 650866 301300 650898
rect 389760 651454 390108 651486
rect 389760 651218 389816 651454
rect 390052 651218 390108 651454
rect 389760 651134 390108 651218
rect 389760 650898 389816 651134
rect 390052 650898 390108 651134
rect 389760 650866 390108 650898
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 300272 619954 300620 619986
rect 300272 619718 300328 619954
rect 300564 619718 300620 619954
rect 300272 619634 300620 619718
rect 300272 619398 300328 619634
rect 300564 619398 300620 619634
rect 300272 619366 300620 619398
rect 390440 619954 390788 619986
rect 390440 619718 390496 619954
rect 390732 619718 390788 619954
rect 390440 619634 390788 619718
rect 390440 619398 390496 619634
rect 390732 619398 390788 619634
rect 390440 619366 390788 619398
rect 300952 615454 301300 615486
rect 300952 615218 301008 615454
rect 301244 615218 301300 615454
rect 300952 615134 301300 615218
rect 300952 614898 301008 615134
rect 301244 614898 301300 615134
rect 300952 614866 301300 614898
rect 389760 615454 390108 615486
rect 389760 615218 389816 615454
rect 390052 615218 390108 615454
rect 389760 615134 390108 615218
rect 389760 614898 389816 615134
rect 390052 614898 390108 615134
rect 389760 614866 390108 614898
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 312928 599450 312988 600100
rect 312862 599390 312988 599450
rect 314288 599450 314348 600100
rect 315376 599450 315436 600100
rect 317688 599586 317748 600100
rect 314288 599390 314394 599450
rect 312862 596597 312922 599390
rect 314334 596869 314394 599390
rect 315254 599390 315436 599450
rect 317646 599526 317748 599586
rect 318912 599586 318972 600100
rect 320000 599586 320060 600100
rect 321088 599586 321148 600100
rect 322312 599586 322372 600100
rect 323400 599586 323460 600100
rect 318912 599526 318994 599586
rect 320000 599526 320098 599586
rect 321088 599526 321202 599586
rect 315254 597005 315314 599390
rect 317646 597549 317706 599526
rect 318934 597549 318994 599526
rect 320038 597549 320098 599526
rect 321142 597549 321202 599526
rect 322246 599526 322372 599586
rect 323350 599526 323460 599586
rect 324760 599586 324820 600100
rect 325304 599586 325364 600100
rect 324760 599526 324882 599586
rect 322246 597549 322306 599526
rect 323350 597549 323410 599526
rect 317643 597548 317709 597549
rect 317643 597484 317644 597548
rect 317708 597484 317709 597548
rect 317643 597483 317709 597484
rect 318931 597548 318997 597549
rect 318931 597484 318932 597548
rect 318996 597484 318997 597548
rect 318931 597483 318997 597484
rect 320035 597548 320101 597549
rect 320035 597484 320036 597548
rect 320100 597484 320101 597548
rect 320035 597483 320101 597484
rect 321139 597548 321205 597549
rect 321139 597484 321140 597548
rect 321204 597484 321205 597548
rect 321139 597483 321205 597484
rect 322243 597548 322309 597549
rect 322243 597484 322244 597548
rect 322308 597484 322309 597548
rect 322243 597483 322309 597484
rect 323347 597548 323413 597549
rect 323347 597484 323348 597548
rect 323412 597484 323413 597548
rect 323347 597483 323413 597484
rect 324822 597413 324882 599526
rect 325190 599526 325364 599586
rect 325712 599586 325772 600100
rect 330472 599586 330532 600100
rect 325712 599526 325802 599586
rect 330472 599526 330586 599586
rect 325190 597549 325250 599526
rect 325742 597549 325802 599526
rect 330526 597549 330586 599526
rect 335504 599450 335564 600100
rect 340536 599450 340596 600100
rect 335126 599390 335564 599450
rect 340462 599390 340596 599450
rect 345568 599450 345628 600100
rect 350464 599450 350524 600100
rect 355496 599450 355556 600100
rect 360528 599450 360588 600100
rect 345568 599390 345674 599450
rect 325187 597548 325253 597549
rect 325187 597484 325188 597548
rect 325252 597484 325253 597548
rect 325187 597483 325253 597484
rect 325739 597548 325805 597549
rect 325739 597484 325740 597548
rect 325804 597484 325805 597548
rect 325739 597483 325805 597484
rect 330523 597548 330589 597549
rect 330523 597484 330524 597548
rect 330588 597484 330589 597548
rect 330523 597483 330589 597484
rect 324819 597412 324885 597413
rect 324819 597348 324820 597412
rect 324884 597348 324885 597412
rect 324819 597347 324885 597348
rect 315251 597004 315317 597005
rect 315251 596940 315252 597004
rect 315316 596940 315317 597004
rect 315251 596939 315317 596940
rect 314331 596868 314397 596869
rect 314331 596804 314332 596868
rect 314396 596804 314397 596868
rect 314331 596803 314397 596804
rect 312859 596596 312925 596597
rect 312859 596532 312860 596596
rect 312924 596532 312925 596596
rect 312859 596531 312925 596532
rect 335126 596325 335186 599390
rect 340462 597005 340522 599390
rect 345614 597549 345674 599390
rect 350398 599390 350524 599450
rect 354446 599390 355556 599450
rect 360518 599390 360588 599450
rect 345611 597548 345677 597549
rect 345611 597484 345612 597548
rect 345676 597484 345677 597548
rect 345611 597483 345677 597484
rect 350398 597141 350458 599390
rect 350395 597140 350461 597141
rect 350395 597076 350396 597140
rect 350460 597076 350461 597140
rect 350395 597075 350461 597076
rect 340459 597004 340525 597005
rect 340459 596940 340460 597004
rect 340524 596940 340525 597004
rect 340459 596939 340525 596940
rect 354446 596325 354506 599390
rect 360518 597549 360578 599390
rect 360515 597548 360581 597549
rect 360515 597484 360516 597548
rect 360580 597484 360581 597548
rect 360515 597483 360581 597484
rect 335123 596324 335189 596325
rect 335123 596260 335124 596324
rect 335188 596260 335189 596324
rect 335123 596259 335189 596260
rect 354443 596324 354509 596325
rect 354443 596260 354444 596324
rect 354508 596260 354509 596324
rect 354443 596259 354509 596260
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 300272 547954 300620 547986
rect 300272 547718 300328 547954
rect 300564 547718 300620 547954
rect 300272 547634 300620 547718
rect 300272 547398 300328 547634
rect 300564 547398 300620 547634
rect 300272 547366 300620 547398
rect 390440 547954 390788 547986
rect 390440 547718 390496 547954
rect 390732 547718 390788 547954
rect 390440 547634 390788 547718
rect 390440 547398 390496 547634
rect 390732 547398 390788 547634
rect 390440 547366 390788 547398
rect 300952 543454 301300 543486
rect 300952 543218 301008 543454
rect 301244 543218 301300 543454
rect 300952 543134 301300 543218
rect 300952 542898 301008 543134
rect 301244 542898 301300 543134
rect 300952 542866 301300 542898
rect 389760 543454 390108 543486
rect 389760 543218 389816 543454
rect 390052 543218 390108 543454
rect 389760 543134 390108 543218
rect 389760 542898 389816 543134
rect 390052 542898 390108 543134
rect 389760 542866 390108 542898
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 300272 511954 300620 511986
rect 300272 511718 300328 511954
rect 300564 511718 300620 511954
rect 300272 511634 300620 511718
rect 300272 511398 300328 511634
rect 300564 511398 300620 511634
rect 300272 511366 300620 511398
rect 390440 511954 390788 511986
rect 390440 511718 390496 511954
rect 390732 511718 390788 511954
rect 390440 511634 390788 511718
rect 390440 511398 390496 511634
rect 390732 511398 390788 511634
rect 390440 511366 390788 511398
rect 300952 507454 301300 507486
rect 300952 507218 301008 507454
rect 301244 507218 301300 507454
rect 300952 507134 301300 507218
rect 300952 506898 301008 507134
rect 301244 506898 301300 507134
rect 300952 506866 301300 506898
rect 389760 507454 390108 507486
rect 389760 507218 389816 507454
rect 390052 507218 390108 507454
rect 389760 507134 390108 507218
rect 389760 506898 389816 507134
rect 390052 506898 390108 507134
rect 389760 506866 390108 506898
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 312928 489930 312988 490106
rect 314288 489930 314348 490106
rect 315376 489930 315436 490106
rect 317688 489930 317748 490106
rect 312928 489870 313106 489930
rect 314288 489870 314394 489930
rect 315376 489870 315498 489930
rect 313046 487933 313106 489870
rect 314334 488477 314394 489870
rect 315438 488477 315498 489870
rect 317646 489870 317748 489930
rect 318912 489930 318972 490106
rect 320000 489930 320060 490106
rect 321088 489930 321148 490106
rect 322312 489930 322372 490106
rect 323400 489930 323460 490106
rect 318912 489870 318994 489930
rect 320000 489870 320098 489930
rect 321088 489870 321202 489930
rect 314331 488476 314397 488477
rect 314331 488412 314332 488476
rect 314396 488412 314397 488476
rect 314331 488411 314397 488412
rect 315435 488476 315501 488477
rect 315435 488412 315436 488476
rect 315500 488412 315501 488476
rect 315435 488411 315501 488412
rect 313043 487932 313109 487933
rect 313043 487868 313044 487932
rect 313108 487868 313109 487932
rect 313043 487867 313109 487868
rect 317646 487253 317706 489870
rect 318934 487389 318994 489870
rect 318931 487388 318997 487389
rect 318931 487324 318932 487388
rect 318996 487324 318997 487388
rect 318931 487323 318997 487324
rect 320038 487253 320098 489870
rect 321142 487525 321202 489870
rect 322246 489870 322372 489930
rect 323350 489870 323460 489930
rect 324760 489930 324820 490106
rect 325304 489930 325364 490106
rect 324760 489870 324882 489930
rect 321139 487524 321205 487525
rect 321139 487460 321140 487524
rect 321204 487460 321205 487524
rect 321139 487459 321205 487460
rect 322246 487253 322306 489870
rect 323350 488477 323410 489870
rect 323347 488476 323413 488477
rect 323347 488412 323348 488476
rect 323412 488412 323413 488476
rect 323347 488411 323413 488412
rect 324822 487525 324882 489870
rect 325190 489870 325364 489930
rect 325712 489930 325772 490106
rect 330472 489930 330532 490106
rect 335504 489930 335564 490106
rect 340536 489930 340596 490106
rect 325712 489870 325802 489930
rect 330472 489870 330586 489930
rect 324819 487524 324885 487525
rect 324819 487460 324820 487524
rect 324884 487460 324885 487524
rect 324819 487459 324885 487460
rect 325190 487253 325250 489870
rect 325742 487253 325802 489870
rect 330526 487253 330586 489870
rect 335494 489870 335564 489930
rect 340462 489870 340596 489930
rect 345568 489930 345628 490106
rect 350464 489930 350524 490106
rect 345568 489870 345674 489930
rect 335494 487253 335554 489870
rect 340462 487253 340522 489870
rect 345614 487253 345674 489870
rect 350398 489870 350524 489930
rect 355496 489930 355556 490106
rect 360528 489930 360588 490106
rect 355496 489870 355610 489930
rect 350398 487253 350458 489870
rect 355550 487253 355610 489870
rect 360518 489870 360588 489930
rect 360518 487253 360578 489870
rect 317643 487252 317709 487253
rect 317643 487188 317644 487252
rect 317708 487188 317709 487252
rect 317643 487187 317709 487188
rect 320035 487252 320101 487253
rect 320035 487188 320036 487252
rect 320100 487188 320101 487252
rect 320035 487187 320101 487188
rect 322243 487252 322309 487253
rect 322243 487188 322244 487252
rect 322308 487188 322309 487252
rect 322243 487187 322309 487188
rect 325187 487252 325253 487253
rect 325187 487188 325188 487252
rect 325252 487188 325253 487252
rect 325187 487187 325253 487188
rect 325739 487252 325805 487253
rect 325739 487188 325740 487252
rect 325804 487188 325805 487252
rect 325739 487187 325805 487188
rect 330523 487252 330589 487253
rect 330523 487188 330524 487252
rect 330588 487188 330589 487252
rect 330523 487187 330589 487188
rect 335491 487252 335557 487253
rect 335491 487188 335492 487252
rect 335556 487188 335557 487252
rect 335491 487187 335557 487188
rect 340459 487252 340525 487253
rect 340459 487188 340460 487252
rect 340524 487188 340525 487252
rect 340459 487187 340525 487188
rect 345611 487252 345677 487253
rect 345611 487188 345612 487252
rect 345676 487188 345677 487252
rect 345611 487187 345677 487188
rect 350395 487252 350461 487253
rect 350395 487188 350396 487252
rect 350460 487188 350461 487252
rect 350395 487187 350461 487188
rect 355547 487252 355613 487253
rect 355547 487188 355548 487252
rect 355612 487188 355613 487252
rect 355547 487187 355613 487188
rect 360515 487252 360581 487253
rect 360515 487188 360516 487252
rect 360580 487188 360581 487252
rect 360515 487187 360581 487188
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 388794 462454 389414 488000
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 382227 454340 382293 454341
rect 382227 454276 382228 454340
rect 382292 454276 382293 454340
rect 382227 454275 382293 454276
rect 378731 454204 378797 454205
rect 378731 454140 378732 454204
rect 378796 454140 378797 454204
rect 378731 454139 378797 454140
rect 378734 453930 378794 454139
rect 379099 454068 379165 454069
rect 379099 454004 379100 454068
rect 379164 454004 379165 454068
rect 379099 454003 379165 454004
rect 379102 453930 379162 454003
rect 378734 453870 379162 453930
rect 298507 446452 298573 446453
rect 298507 446388 298508 446452
rect 298572 446388 298573 446452
rect 298507 446387 298573 446388
rect 295931 444412 295997 444413
rect 295931 444348 295932 444412
rect 295996 444348 295997 444412
rect 295931 444347 295997 444348
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 295934 19413 295994 444347
rect 295931 19412 295997 19413
rect 295931 19348 295932 19412
rect 295996 19348 295997 19412
rect 295931 19347 295997 19348
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 298510 5677 298570 446387
rect 382230 441630 382290 454275
rect 382230 441570 383394 441630
rect 319568 439954 319888 439986
rect 319568 439718 319610 439954
rect 319846 439718 319888 439954
rect 319568 439634 319888 439718
rect 319568 439398 319610 439634
rect 319846 439398 319888 439634
rect 319568 439366 319888 439398
rect 350288 439954 350608 439986
rect 350288 439718 350330 439954
rect 350566 439718 350608 439954
rect 350288 439634 350608 439718
rect 350288 439398 350330 439634
rect 350566 439398 350608 439634
rect 350288 439366 350608 439398
rect 381008 439954 381328 439986
rect 381008 439718 381050 439954
rect 381286 439718 381328 439954
rect 381008 439634 381328 439718
rect 381008 439398 381050 439634
rect 381286 439398 381328 439634
rect 381008 439366 381328 439398
rect 304208 435454 304528 435486
rect 304208 435218 304250 435454
rect 304486 435218 304528 435454
rect 304208 435134 304528 435218
rect 304208 434898 304250 435134
rect 304486 434898 304528 435134
rect 304208 434866 304528 434898
rect 334928 435454 335248 435486
rect 334928 435218 334970 435454
rect 335206 435218 335248 435454
rect 334928 435134 335248 435218
rect 334928 434898 334970 435134
rect 335206 434898 335248 435134
rect 334928 434866 335248 434898
rect 365648 435454 365968 435486
rect 365648 435218 365690 435454
rect 365926 435218 365968 435454
rect 365648 435134 365968 435218
rect 365648 434898 365690 435134
rect 365926 434898 365968 435134
rect 365648 434866 365968 434898
rect 383334 425781 383394 441570
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 383331 425780 383397 425781
rect 383331 425716 383332 425780
rect 383396 425716 383397 425780
rect 383331 425715 383397 425716
rect 319568 403954 319888 403986
rect 319568 403718 319610 403954
rect 319846 403718 319888 403954
rect 319568 403634 319888 403718
rect 319568 403398 319610 403634
rect 319846 403398 319888 403634
rect 319568 403366 319888 403398
rect 350288 403954 350608 403986
rect 350288 403718 350330 403954
rect 350566 403718 350608 403954
rect 350288 403634 350608 403718
rect 350288 403398 350330 403634
rect 350566 403398 350608 403634
rect 350288 403366 350608 403398
rect 381008 403954 381328 403986
rect 381008 403718 381050 403954
rect 381286 403718 381328 403954
rect 381008 403634 381328 403718
rect 381008 403398 381050 403634
rect 381286 403398 381328 403634
rect 381008 403366 381328 403398
rect 332547 401028 332613 401029
rect 332547 400964 332548 401028
rect 332612 400964 332613 401028
rect 332547 400963 332613 400964
rect 332550 400621 332610 400963
rect 332547 400620 332613 400621
rect 332547 400556 332548 400620
rect 332612 400556 332613 400620
rect 332547 400555 332613 400556
rect 298794 372454 299414 398000
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 5676 298573 5677
rect 298507 5612 298508 5676
rect 298572 5612 298573 5676
rect 298507 5611 298573 5612
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 376954 303914 398000
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 381454 308414 398000
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 385954 312914 398000
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 390454 317414 398000
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 394954 321914 398000
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 367954 330914 398000
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 372454 335414 398000
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 376954 339914 398000
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 385954 348914 398000
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 390454 353414 398000
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 394954 357914 398000
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 363454 362414 398000
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 367954 366914 398000
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 372454 371414 398000
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 376954 375914 398000
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 381454 380414 398000
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 385954 384914 398000
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 691292 411914 700398
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 691292 438914 691398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 691292 443414 695898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 691292 447914 700398
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 691292 474914 691398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 691292 479414 695898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 691292 483914 700398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 410952 687454 411300 687486
rect 410952 687218 411008 687454
rect 411244 687218 411300 687454
rect 410952 687134 411300 687218
rect 410952 686898 411008 687134
rect 411244 686898 411300 687134
rect 410952 686866 411300 686898
rect 499760 687454 500108 687486
rect 499760 687218 499816 687454
rect 500052 687218 500108 687454
rect 499760 687134 500108 687218
rect 499760 686898 499816 687134
rect 500052 686898 500108 687134
rect 499760 686866 500108 686898
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 410272 655954 410620 655986
rect 410272 655718 410328 655954
rect 410564 655718 410620 655954
rect 410272 655634 410620 655718
rect 410272 655398 410328 655634
rect 410564 655398 410620 655634
rect 410272 655366 410620 655398
rect 500440 655954 500788 655986
rect 500440 655718 500496 655954
rect 500732 655718 500788 655954
rect 500440 655634 500788 655718
rect 500440 655398 500496 655634
rect 500732 655398 500788 655634
rect 500440 655366 500788 655398
rect 410952 651454 411300 651486
rect 410952 651218 411008 651454
rect 411244 651218 411300 651454
rect 410952 651134 411300 651218
rect 410952 650898 411008 651134
rect 411244 650898 411300 651134
rect 410952 650866 411300 650898
rect 499760 651454 500108 651486
rect 499760 651218 499816 651454
rect 500052 651218 500108 651454
rect 499760 651134 500108 651218
rect 499760 650898 499816 651134
rect 500052 650898 500108 651134
rect 499760 650866 500108 650898
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 410272 619954 410620 619986
rect 410272 619718 410328 619954
rect 410564 619718 410620 619954
rect 410272 619634 410620 619718
rect 410272 619398 410328 619634
rect 410564 619398 410620 619634
rect 410272 619366 410620 619398
rect 500440 619954 500788 619986
rect 500440 619718 500496 619954
rect 500732 619718 500788 619954
rect 500440 619634 500788 619718
rect 500440 619398 500496 619634
rect 500732 619398 500788 619634
rect 500440 619366 500788 619398
rect 410952 615454 411300 615486
rect 410952 615218 411008 615454
rect 411244 615218 411300 615454
rect 410952 615134 411300 615218
rect 410952 614898 411008 615134
rect 411244 614898 411300 615134
rect 410952 614866 411300 614898
rect 499760 615454 500108 615486
rect 499760 615218 499816 615454
rect 500052 615218 500108 615454
rect 499760 615134 500108 615218
rect 499760 614898 499816 615134
rect 500052 614898 500108 615134
rect 499760 614866 500108 614898
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 422928 599450 422988 600100
rect 424288 599450 424348 600100
rect 425376 599450 425436 600100
rect 427688 599450 427748 600100
rect 422894 599390 422988 599450
rect 424182 599390 424348 599450
rect 425286 599390 425436 599450
rect 427678 599390 427748 599450
rect 428912 599450 428972 600100
rect 430000 599450 430060 600100
rect 431088 599450 431148 600100
rect 432312 599450 432372 600100
rect 433400 599450 433460 600100
rect 434760 599450 434820 600100
rect 435304 599450 435364 600100
rect 435712 599450 435772 600100
rect 440472 599450 440532 600100
rect 428912 599390 429026 599450
rect 422894 597277 422954 599390
rect 422891 597276 422957 597277
rect 422891 597212 422892 597276
rect 422956 597212 422957 597276
rect 422891 597211 422957 597212
rect 424182 597005 424242 599390
rect 424179 597004 424245 597005
rect 424179 596940 424180 597004
rect 424244 596940 424245 597004
rect 424179 596939 424245 596940
rect 425286 596461 425346 599390
rect 427678 597277 427738 599390
rect 428966 597277 429026 599390
rect 429886 599390 430060 599450
rect 430990 599390 431148 599450
rect 431726 599390 432372 599450
rect 433382 599390 433460 599450
rect 434670 599390 434820 599450
rect 435222 599390 435364 599450
rect 435590 599390 435772 599450
rect 440374 599390 440532 599450
rect 445504 599450 445564 600100
rect 450536 599450 450596 600100
rect 455568 599450 455628 600100
rect 460464 599450 460524 600100
rect 465496 599450 465556 600100
rect 470528 599450 470588 600100
rect 445504 599390 445586 599450
rect 427675 597276 427741 597277
rect 427675 597212 427676 597276
rect 427740 597212 427741 597276
rect 427675 597211 427741 597212
rect 428963 597276 429029 597277
rect 428963 597212 428964 597276
rect 429028 597212 429029 597276
rect 428963 597211 429029 597212
rect 429886 597141 429946 599390
rect 430990 597277 431050 599390
rect 430987 597276 431053 597277
rect 430987 597212 430988 597276
rect 431052 597212 431053 597276
rect 430987 597211 431053 597212
rect 429883 597140 429949 597141
rect 429883 597076 429884 597140
rect 429948 597076 429949 597140
rect 429883 597075 429949 597076
rect 431726 597005 431786 599390
rect 433382 597005 433442 599390
rect 434670 597005 434730 599390
rect 431723 597004 431789 597005
rect 431723 596940 431724 597004
rect 431788 596940 431789 597004
rect 431723 596939 431789 596940
rect 433379 597004 433445 597005
rect 433379 596940 433380 597004
rect 433444 596940 433445 597004
rect 433379 596939 433445 596940
rect 434667 597004 434733 597005
rect 434667 596940 434668 597004
rect 434732 596940 434733 597004
rect 434667 596939 434733 596940
rect 435222 596733 435282 599390
rect 435590 597413 435650 599390
rect 440374 597549 440434 599390
rect 440371 597548 440437 597549
rect 440371 597484 440372 597548
rect 440436 597484 440437 597548
rect 440371 597483 440437 597484
rect 435587 597412 435653 597413
rect 435587 597348 435588 597412
rect 435652 597348 435653 597412
rect 435587 597347 435653 597348
rect 445526 596733 445586 599390
rect 450494 599390 450596 599450
rect 455462 599390 455628 599450
rect 460430 599390 460524 599450
rect 465398 599390 465556 599450
rect 470366 599390 470588 599450
rect 450494 597549 450554 599390
rect 450491 597548 450557 597549
rect 450491 597484 450492 597548
rect 450556 597484 450557 597548
rect 450491 597483 450557 597484
rect 435219 596732 435285 596733
rect 435219 596668 435220 596732
rect 435284 596668 435285 596732
rect 435219 596667 435285 596668
rect 445523 596732 445589 596733
rect 445523 596668 445524 596732
rect 445588 596668 445589 596732
rect 445523 596667 445589 596668
rect 425283 596460 425349 596461
rect 425283 596396 425284 596460
rect 425348 596396 425349 596460
rect 425283 596395 425349 596396
rect 455462 596325 455522 599390
rect 460430 597549 460490 599390
rect 460427 597548 460493 597549
rect 460427 597484 460428 597548
rect 460492 597484 460493 597548
rect 460427 597483 460493 597484
rect 465398 596869 465458 599390
rect 465395 596868 465461 596869
rect 465395 596804 465396 596868
rect 465460 596804 465461 596868
rect 465395 596803 465461 596804
rect 470366 596325 470426 599390
rect 455459 596324 455525 596325
rect 455459 596260 455460 596324
rect 455524 596260 455525 596324
rect 455459 596259 455525 596260
rect 470363 596324 470429 596325
rect 470363 596260 470364 596324
rect 470428 596260 470429 596324
rect 470363 596259 470429 596260
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 410272 547954 410620 547986
rect 410272 547718 410328 547954
rect 410564 547718 410620 547954
rect 410272 547634 410620 547718
rect 410272 547398 410328 547634
rect 410564 547398 410620 547634
rect 410272 547366 410620 547398
rect 500440 547954 500788 547986
rect 500440 547718 500496 547954
rect 500732 547718 500788 547954
rect 500440 547634 500788 547718
rect 500440 547398 500496 547634
rect 500732 547398 500788 547634
rect 500440 547366 500788 547398
rect 410952 543454 411300 543486
rect 410952 543218 411008 543454
rect 411244 543218 411300 543454
rect 410952 543134 411300 543218
rect 410952 542898 411008 543134
rect 411244 542898 411300 543134
rect 410952 542866 411300 542898
rect 499760 543454 500108 543486
rect 499760 543218 499816 543454
rect 500052 543218 500108 543454
rect 499760 543134 500108 543218
rect 499760 542898 499816 543134
rect 500052 542898 500108 543134
rect 499760 542866 500108 542898
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 407803 526692 407869 526693
rect 407803 526628 407804 526692
rect 407868 526628 407869 526692
rect 407803 526627 407869 526628
rect 407619 523700 407685 523701
rect 407619 523636 407620 523700
rect 407684 523636 407685 523700
rect 407619 523635 407685 523636
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 407622 489837 407682 523635
rect 407619 489836 407685 489837
rect 407619 489772 407620 489836
rect 407684 489772 407685 489836
rect 407619 489771 407685 489772
rect 407806 488069 407866 526627
rect 410272 511954 410620 511986
rect 410272 511718 410328 511954
rect 410564 511718 410620 511954
rect 410272 511634 410620 511718
rect 410272 511398 410328 511634
rect 410564 511398 410620 511634
rect 410272 511366 410620 511398
rect 500440 511954 500788 511986
rect 500440 511718 500496 511954
rect 500732 511718 500788 511954
rect 500440 511634 500788 511718
rect 500440 511398 500496 511634
rect 500732 511398 500788 511634
rect 500440 511366 500788 511398
rect 410952 507454 411300 507486
rect 410952 507218 411008 507454
rect 411244 507218 411300 507454
rect 410952 507134 411300 507218
rect 410952 506898 411008 507134
rect 411244 506898 411300 507134
rect 410952 506866 411300 506898
rect 499760 507454 500108 507486
rect 499760 507218 499816 507454
rect 500052 507218 500108 507454
rect 499760 507134 500108 507218
rect 499760 506898 499816 507134
rect 500052 506898 500108 507134
rect 499760 506866 500108 506898
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 422928 489930 422988 490106
rect 424288 489930 424348 490106
rect 425376 489930 425436 490106
rect 427688 489930 427748 490106
rect 422894 489870 422988 489930
rect 424182 489870 424348 489930
rect 425286 489870 425436 489930
rect 427678 489870 427748 489930
rect 428912 489930 428972 490106
rect 430000 489930 430060 490106
rect 431088 489930 431148 490106
rect 432312 489930 432372 490106
rect 433400 489930 433460 490106
rect 428912 489870 429026 489930
rect 422894 488477 422954 489870
rect 424182 488477 424242 489870
rect 425286 488477 425346 489870
rect 422891 488476 422957 488477
rect 422891 488412 422892 488476
rect 422956 488412 422957 488476
rect 422891 488411 422957 488412
rect 424179 488476 424245 488477
rect 424179 488412 424180 488476
rect 424244 488412 424245 488476
rect 424179 488411 424245 488412
rect 425283 488476 425349 488477
rect 425283 488412 425284 488476
rect 425348 488412 425349 488476
rect 425283 488411 425349 488412
rect 407803 488068 407869 488069
rect 407803 488004 407804 488068
rect 407868 488004 407869 488068
rect 407803 488003 407869 488004
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 484954 411914 488000
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 453454 416414 488000
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 457954 420914 488000
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 462454 425414 488000
rect 427678 487661 427738 489870
rect 428966 487797 429026 489870
rect 429886 489870 430060 489930
rect 430990 489870 431148 489930
rect 432278 489870 432372 489930
rect 433382 489870 433460 489930
rect 434760 489930 434820 490106
rect 435304 489930 435364 490106
rect 435712 489930 435772 490106
rect 440472 489930 440532 490106
rect 434760 489870 434914 489930
rect 429886 488205 429946 489870
rect 429883 488204 429949 488205
rect 429883 488140 429884 488204
rect 429948 488140 429949 488204
rect 429883 488139 429949 488140
rect 428963 487796 429029 487797
rect 428963 487732 428964 487796
rect 429028 487732 429029 487796
rect 428963 487731 429029 487732
rect 427675 487660 427741 487661
rect 427675 487596 427676 487660
rect 427740 487596 427741 487660
rect 427675 487595 427741 487596
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 466954 429914 488000
rect 430990 487525 431050 489870
rect 432278 487525 432338 489870
rect 433382 487525 433442 489870
rect 430987 487524 431053 487525
rect 430987 487460 430988 487524
rect 431052 487460 431053 487524
rect 430987 487459 431053 487460
rect 432275 487524 432341 487525
rect 432275 487460 432276 487524
rect 432340 487460 432341 487524
rect 432275 487459 432341 487460
rect 433379 487524 433445 487525
rect 433379 487460 433380 487524
rect 433444 487460 433445 487524
rect 433379 487459 433445 487460
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 471454 434414 488000
rect 434854 487525 434914 489870
rect 435222 489870 435364 489930
rect 435590 489870 435772 489930
rect 440374 489870 440532 489930
rect 445504 489930 445564 490106
rect 450536 489930 450596 490106
rect 455568 489930 455628 490106
rect 460464 489930 460524 490106
rect 465496 489930 465556 490106
rect 445504 489870 445586 489930
rect 434851 487524 434917 487525
rect 434851 487460 434852 487524
rect 434916 487460 434917 487524
rect 434851 487459 434917 487460
rect 435222 487253 435282 489870
rect 435590 487661 435650 489870
rect 435587 487660 435653 487661
rect 435587 487596 435588 487660
rect 435652 487596 435653 487660
rect 435587 487595 435653 487596
rect 435219 487252 435285 487253
rect 435219 487188 435220 487252
rect 435284 487188 435285 487252
rect 435219 487187 435285 487188
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 475954 438914 488000
rect 440374 487253 440434 489870
rect 440371 487252 440437 487253
rect 440371 487188 440372 487252
rect 440436 487188 440437 487252
rect 440371 487187 440437 487188
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 480454 443414 488000
rect 445526 487253 445586 489870
rect 450494 489870 450596 489930
rect 455462 489870 455628 489930
rect 460430 489870 460524 489930
rect 465398 489870 465556 489930
rect 470528 489930 470588 490106
rect 470528 489870 470794 489930
rect 445523 487252 445589 487253
rect 445523 487188 445524 487252
rect 445588 487188 445589 487252
rect 445523 487187 445589 487188
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 484954 447914 488000
rect 450494 487253 450554 489870
rect 450491 487252 450557 487253
rect 450491 487188 450492 487252
rect 450556 487188 450557 487252
rect 450491 487187 450557 487188
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 453454 452414 488000
rect 455462 487253 455522 489870
rect 455459 487252 455525 487253
rect 455459 487188 455460 487252
rect 455524 487188 455525 487252
rect 455459 487187 455525 487188
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 457954 456914 488000
rect 460430 487253 460490 489870
rect 465398 488341 465458 489870
rect 465395 488340 465461 488341
rect 465395 488276 465396 488340
rect 465460 488276 465461 488340
rect 465395 488275 465461 488276
rect 460427 487252 460493 487253
rect 460427 487188 460428 487252
rect 460492 487188 460493 487252
rect 460427 487187 460493 487188
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 462454 461414 488000
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 466954 465914 488000
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 471454 470414 488000
rect 470734 487253 470794 489870
rect 470731 487252 470797 487253
rect 470731 487188 470732 487252
rect 470796 487188 470797 487252
rect 470731 487187 470797 487188
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 475954 474914 488000
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 480454 479414 488000
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 484954 483914 488000
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 453454 488414 488000
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 457954 492914 488000
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 462454 497414 488000
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 466954 501914 488000
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 81008 687218 81244 687454
rect 81008 686898 81244 687134
rect 169816 687218 170052 687454
rect 169816 686898 170052 687134
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 80328 655718 80564 655954
rect 80328 655398 80564 655634
rect 170496 655718 170732 655954
rect 170496 655398 170732 655634
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 81008 651218 81244 651454
rect 81008 650898 81244 651134
rect 169816 651218 170052 651454
rect 169816 650898 170052 651134
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 80328 619718 80564 619954
rect 80328 619398 80564 619634
rect 170496 619718 170732 619954
rect 170496 619398 170732 619634
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 81008 615218 81244 615454
rect 81008 614898 81244 615134
rect 169816 615218 170052 615454
rect 169816 614898 170052 615134
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 80328 547718 80564 547954
rect 80328 547398 80564 547634
rect 170496 547718 170732 547954
rect 170496 547398 170732 547634
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 81008 543218 81244 543454
rect 81008 542898 81244 543134
rect 169816 543218 170052 543454
rect 169816 542898 170052 543134
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 80328 511718 80564 511954
rect 80328 511398 80564 511634
rect 170496 511718 170732 511954
rect 170496 511398 170732 511634
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 81008 507218 81244 507454
rect 81008 506898 81244 507134
rect 169816 507218 170052 507454
rect 169816 506898 170052 507134
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 191008 687218 191244 687454
rect 191008 686898 191244 687134
rect 279816 687218 280052 687454
rect 279816 686898 280052 687134
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 190328 655718 190564 655954
rect 190328 655398 190564 655634
rect 280496 655718 280732 655954
rect 280496 655398 280732 655634
rect 191008 651218 191244 651454
rect 191008 650898 191244 651134
rect 279816 651218 280052 651454
rect 279816 650898 280052 651134
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 190328 619718 190564 619954
rect 190328 619398 190564 619634
rect 280496 619718 280732 619954
rect 280496 619398 280732 619634
rect 191008 615218 191244 615454
rect 191008 614898 191244 615134
rect 279816 615218 280052 615454
rect 279816 614898 280052 615134
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 190328 547718 190564 547954
rect 190328 547398 190564 547634
rect 280496 547718 280732 547954
rect 280496 547398 280732 547634
rect 191008 543218 191244 543454
rect 191008 542898 191244 543134
rect 279816 543218 280052 543454
rect 279816 542898 280052 543134
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 190328 511718 190564 511954
rect 190328 511398 190564 511634
rect 280496 511718 280732 511954
rect 280496 511398 280732 511634
rect 191008 507218 191244 507454
rect 191008 506898 191244 507134
rect 279816 507218 280052 507454
rect 279816 506898 280052 507134
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 219610 439718 219846 439954
rect 219610 439398 219846 439634
rect 250330 439718 250566 439954
rect 250330 439398 250566 439634
rect 204250 435218 204486 435454
rect 204250 434898 204486 435134
rect 234970 435218 235206 435454
rect 234970 434898 235206 435134
rect 219610 403718 219846 403954
rect 219610 403398 219846 403634
rect 250330 403718 250566 403954
rect 250330 403398 250566 403634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 301008 687218 301244 687454
rect 301008 686898 301244 687134
rect 389816 687218 390052 687454
rect 389816 686898 390052 687134
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 300328 655718 300564 655954
rect 300328 655398 300564 655634
rect 390496 655718 390732 655954
rect 390496 655398 390732 655634
rect 301008 651218 301244 651454
rect 301008 650898 301244 651134
rect 389816 651218 390052 651454
rect 389816 650898 390052 651134
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 300328 619718 300564 619954
rect 300328 619398 300564 619634
rect 390496 619718 390732 619954
rect 390496 619398 390732 619634
rect 301008 615218 301244 615454
rect 301008 614898 301244 615134
rect 389816 615218 390052 615454
rect 389816 614898 390052 615134
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 300328 547718 300564 547954
rect 300328 547398 300564 547634
rect 390496 547718 390732 547954
rect 390496 547398 390732 547634
rect 301008 543218 301244 543454
rect 301008 542898 301244 543134
rect 389816 543218 390052 543454
rect 389816 542898 390052 543134
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 300328 511718 300564 511954
rect 300328 511398 300564 511634
rect 390496 511718 390732 511954
rect 390496 511398 390732 511634
rect 301008 507218 301244 507454
rect 301008 506898 301244 507134
rect 389816 507218 390052 507454
rect 389816 506898 390052 507134
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 319610 439718 319846 439954
rect 319610 439398 319846 439634
rect 350330 439718 350566 439954
rect 350330 439398 350566 439634
rect 381050 439718 381286 439954
rect 381050 439398 381286 439634
rect 304250 435218 304486 435454
rect 304250 434898 304486 435134
rect 334970 435218 335206 435454
rect 334970 434898 335206 435134
rect 365690 435218 365926 435454
rect 365690 434898 365926 435134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 319610 403718 319846 403954
rect 319610 403398 319846 403634
rect 350330 403718 350566 403954
rect 350330 403398 350566 403634
rect 381050 403718 381286 403954
rect 381050 403398 381286 403634
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 411008 687218 411244 687454
rect 411008 686898 411244 687134
rect 499816 687218 500052 687454
rect 499816 686898 500052 687134
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 410328 655718 410564 655954
rect 410328 655398 410564 655634
rect 500496 655718 500732 655954
rect 500496 655398 500732 655634
rect 411008 651218 411244 651454
rect 411008 650898 411244 651134
rect 499816 651218 500052 651454
rect 499816 650898 500052 651134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 410328 619718 410564 619954
rect 410328 619398 410564 619634
rect 500496 619718 500732 619954
rect 500496 619398 500732 619634
rect 411008 615218 411244 615454
rect 411008 614898 411244 615134
rect 499816 615218 500052 615454
rect 499816 614898 500052 615134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 410328 547718 410564 547954
rect 410328 547398 410564 547634
rect 500496 547718 500732 547954
rect 500496 547398 500732 547634
rect 411008 543218 411244 543454
rect 411008 542898 411244 543134
rect 499816 543218 500052 543454
rect 499816 542898 500052 543134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 410328 511718 410564 511954
rect 410328 511398 410564 511634
rect 500496 511718 500732 511954
rect 500496 511398 500732 511634
rect 411008 507218 411244 507454
rect 411008 506898 411244 507134
rect 499816 507218 500052 507454
rect 499816 506898 500052 507134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 81008 687454
rect 81244 687218 169816 687454
rect 170052 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 191008 687454
rect 191244 687218 279816 687454
rect 280052 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 301008 687454
rect 301244 687218 389816 687454
rect 390052 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 411008 687454
rect 411244 687218 499816 687454
rect 500052 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 81008 687134
rect 81244 686898 169816 687134
rect 170052 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 191008 687134
rect 191244 686898 279816 687134
rect 280052 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 301008 687134
rect 301244 686898 389816 687134
rect 390052 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 411008 687134
rect 411244 686898 499816 687134
rect 500052 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 80328 655954
rect 80564 655718 170496 655954
rect 170732 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 190328 655954
rect 190564 655718 280496 655954
rect 280732 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 300328 655954
rect 300564 655718 390496 655954
rect 390732 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 410328 655954
rect 410564 655718 500496 655954
rect 500732 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 80328 655634
rect 80564 655398 170496 655634
rect 170732 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 190328 655634
rect 190564 655398 280496 655634
rect 280732 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 300328 655634
rect 300564 655398 390496 655634
rect 390732 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 410328 655634
rect 410564 655398 500496 655634
rect 500732 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 81008 651454
rect 81244 651218 169816 651454
rect 170052 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 191008 651454
rect 191244 651218 279816 651454
rect 280052 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 301008 651454
rect 301244 651218 389816 651454
rect 390052 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 411008 651454
rect 411244 651218 499816 651454
rect 500052 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 81008 651134
rect 81244 650898 169816 651134
rect 170052 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 191008 651134
rect 191244 650898 279816 651134
rect 280052 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 301008 651134
rect 301244 650898 389816 651134
rect 390052 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 411008 651134
rect 411244 650898 499816 651134
rect 500052 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 80328 619954
rect 80564 619718 170496 619954
rect 170732 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 190328 619954
rect 190564 619718 280496 619954
rect 280732 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 300328 619954
rect 300564 619718 390496 619954
rect 390732 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 410328 619954
rect 410564 619718 500496 619954
rect 500732 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 80328 619634
rect 80564 619398 170496 619634
rect 170732 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 190328 619634
rect 190564 619398 280496 619634
rect 280732 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 300328 619634
rect 300564 619398 390496 619634
rect 390732 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 410328 619634
rect 410564 619398 500496 619634
rect 500732 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 81008 615454
rect 81244 615218 169816 615454
rect 170052 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 191008 615454
rect 191244 615218 279816 615454
rect 280052 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 301008 615454
rect 301244 615218 389816 615454
rect 390052 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 411008 615454
rect 411244 615218 499816 615454
rect 500052 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 81008 615134
rect 81244 614898 169816 615134
rect 170052 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 191008 615134
rect 191244 614898 279816 615134
rect 280052 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 301008 615134
rect 301244 614898 389816 615134
rect 390052 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 411008 615134
rect 411244 614898 499816 615134
rect 500052 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 80328 547954
rect 80564 547718 170496 547954
rect 170732 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 190328 547954
rect 190564 547718 280496 547954
rect 280732 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 300328 547954
rect 300564 547718 390496 547954
rect 390732 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 410328 547954
rect 410564 547718 500496 547954
rect 500732 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 80328 547634
rect 80564 547398 170496 547634
rect 170732 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 190328 547634
rect 190564 547398 280496 547634
rect 280732 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 300328 547634
rect 300564 547398 390496 547634
rect 390732 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 410328 547634
rect 410564 547398 500496 547634
rect 500732 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 81008 543454
rect 81244 543218 169816 543454
rect 170052 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 191008 543454
rect 191244 543218 279816 543454
rect 280052 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 301008 543454
rect 301244 543218 389816 543454
rect 390052 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 411008 543454
rect 411244 543218 499816 543454
rect 500052 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 81008 543134
rect 81244 542898 169816 543134
rect 170052 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 191008 543134
rect 191244 542898 279816 543134
rect 280052 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 301008 543134
rect 301244 542898 389816 543134
rect 390052 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 411008 543134
rect 411244 542898 499816 543134
rect 500052 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 80328 511954
rect 80564 511718 170496 511954
rect 170732 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 190328 511954
rect 190564 511718 280496 511954
rect 280732 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 300328 511954
rect 300564 511718 390496 511954
rect 390732 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 410328 511954
rect 410564 511718 500496 511954
rect 500732 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 80328 511634
rect 80564 511398 170496 511634
rect 170732 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 190328 511634
rect 190564 511398 280496 511634
rect 280732 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 300328 511634
rect 300564 511398 390496 511634
rect 390732 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 410328 511634
rect 410564 511398 500496 511634
rect 500732 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 81008 507454
rect 81244 507218 169816 507454
rect 170052 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 191008 507454
rect 191244 507218 279816 507454
rect 280052 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 301008 507454
rect 301244 507218 389816 507454
rect 390052 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 411008 507454
rect 411244 507218 499816 507454
rect 500052 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 81008 507134
rect 81244 506898 169816 507134
rect 170052 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 191008 507134
rect 191244 506898 279816 507134
rect 280052 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 301008 507134
rect 301244 506898 389816 507134
rect 390052 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 411008 507134
rect 411244 506898 499816 507134
rect 500052 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 219610 439954
rect 219846 439718 250330 439954
rect 250566 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 319610 439954
rect 319846 439718 350330 439954
rect 350566 439718 381050 439954
rect 381286 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 219610 439634
rect 219846 439398 250330 439634
rect 250566 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 319610 439634
rect 319846 439398 350330 439634
rect 350566 439398 381050 439634
rect 381286 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 204250 435454
rect 204486 435218 234970 435454
rect 235206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 304250 435454
rect 304486 435218 334970 435454
rect 335206 435218 365690 435454
rect 365926 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 204250 435134
rect 204486 434898 234970 435134
rect 235206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 304250 435134
rect 304486 434898 334970 435134
rect 335206 434898 365690 435134
rect 365926 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 219610 403954
rect 219846 403718 250330 403954
rect 250566 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 319610 403954
rect 319846 403718 350330 403954
rect 350566 403718 381050 403954
rect 381286 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 219610 403634
rect 219846 403398 250330 403634
rect 250566 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 319610 403634
rect 319846 403398 350330 403634
rect 350566 403398 381050 403634
rect 381286 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use cpu  cpu0
timestamp 0
transform 1 0 300000 0 1 400000
box 0 0 84000 56000
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword0
timestamp 0
transform 1 0 80000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword1
timestamp 0
transform 1 0 190000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword2
timestamp 0
transform 1 0 300000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memHword3
timestamp 0
transform 1 0 410000 0 1 600000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword0
timestamp 0
transform 1 0 80000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword1
timestamp 0
transform 1 0 190000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword2
timestamp 0
transform 1 0 300000 0 1 490000
box 0 0 91060 89292
use sky130_sram_1kbyte_1rw1r_8x1024_8  memLword3
timestamp 0
transform 1 0 410000 0 1 490000
box 0 0 91060 89292
use soc_config  mprj
timestamp 0
transform 1 0 200000 0 1 400000
box 1066 0 64898 44000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 398000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 488000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 691292 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 691292 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 691292 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 691292 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 691292 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 691292 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 691292 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 691292 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 398000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 691292 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 691292 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 488000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 691292 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 398000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 488000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 398000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 488000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 398000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 488000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 398000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 488000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 691292 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 691292 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 691292 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 691292 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 691292 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 691292 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 398000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 691292 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 691292 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 488000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 691292 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 691292 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 691292 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 691292 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 691292 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 446000 231914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 691292 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 446000 267914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 691292 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 691292 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 691292 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 398000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 691292 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 691292 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 691292 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 488000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 691292 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
